VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "|" ;

PROPERTYDEFINITIONS
END PROPERTYDEFINITIONS


MACRO fake_macro_newblue1_o330073
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 1.365 7.315 1.435 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330073

MACRO fake_macro_newblue1_o330074
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 1.365 7.315 1.435 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330074

MACRO fake_macro_newblue1_o330075
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 1.365 7.315 1.435 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330075

MACRO fake_macro_newblue1_o330076
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.765 11.725 72.835 11.795 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330076

MACRO fake_macro_newblue1_o330077
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.765 11.725 72.835 11.795 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330077

MACRO fake_macro_newblue1_o330078
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.765 11.725 72.835 11.795 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330078

MACRO fake_macro_newblue1_o330079
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.045 0.035 73.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 73.045 7.315 73.115 ;
        END
    END p2
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330079

MACRO fake_macro_newblue1_o330080
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.045 0.035 73.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 73.045 7.315 73.115 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p2
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330080

MACRO fake_macro_newblue1_o330081
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330081

MACRO fake_macro_newblue1_o330082
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.045 0.035 73.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 73.045 7.315 73.115 ;
        END
    END p2
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330082

MACRO fake_macro_newblue1_o330085
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330085

MACRO fake_macro_newblue1_o330086
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330086

MACRO fake_macro_newblue1_o330087
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330087

MACRO fake_macro_newblue1_o330088
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330088

MACRO fake_macro_newblue1_o330089
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330089

MACRO fake_macro_newblue1_o330090
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330090

MACRO fake_macro_newblue1_o330091
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330091

MACRO fake_macro_newblue1_o330092
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330092

MACRO fake_macro_newblue1_o330093
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330093

MACRO fake_macro_newblue1_o330094
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330094

MACRO fake_macro_newblue1_o330095
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330095

MACRO fake_macro_newblue1_o330096
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 2.485 3.395 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 2.485 6.755 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 10.045 5.075 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330096

MACRO fake_macro_newblue1_o330097
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 2.485 3.395 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 2.485 6.755 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 10.045 5.075 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330097

MACRO fake_macro_newblue1_o330098
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 2.485 3.395 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 2.485 6.755 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 10.045 5.075 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330098

MACRO fake_macro_newblue1_o330099
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 2.485 3.395 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 2.485 6.755 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 10.045 5.075 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330099

MACRO fake_macro_newblue1_o330100
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 2.485 3.395 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 2.485 6.755 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 10.045 5.075 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330100

MACRO fake_macro_newblue1_o330101
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 2.485 3.395 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 2.485 6.755 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 2.485 11.795 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 10.045 5.075 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330101

MACRO fake_macro_newblue1_o330102
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330102

MACRO fake_macro_newblue1_o330103
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 13.125 7.315 13.195 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330103

MACRO fake_macro_newblue1_o330104
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 13.125 7.315 13.195 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330104

MACRO fake_macro_newblue1_o330105
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 13.125 7.315 13.195 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330105

MACRO fake_macro_newblue1_o330106
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 13.125 7.315 13.195 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330106

MACRO fake_macro_newblue1_o330107
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.765 11.445 72.835 11.515 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.205 73.395 2.275 ;
        END
    END p3
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330107

MACRO fake_macro_newblue1_o330108
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 8.365 2.275 8.435 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330108

MACRO fake_macro_newblue1_o330109
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.485 0.595 2.555 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330109

MACRO fake_macro_newblue1_o330110
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 9.765 10.115 9.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 6.965 7.315 7.035 ;
        END
    END p2
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330110

MACRO fake_macro_newblue1_o330111
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 73.045 6.755 73.115 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 70.245 9.555 70.315 ;
        END
    END p2
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330111

MACRO fake_macro_newblue1_o330112
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 8.925 3.395 8.995 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330112

MACRO fake_macro_newblue1_o330113
    CLASS BLOCK ;
    SIZE 80.64 BY 26.88 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 18.165 2.275 18.235 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 2.485 8.995 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.605 2.275 17.675 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 15.925 2.275 15.995 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.925 2.275 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 10.325 2.275 10.395 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 15.085 2.275 15.155 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 15.645 2.275 15.715 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 0.245 6.755 0.315 ;
        END
    END p9
    PIN p10
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.645 51.555 1.715 ;
        END
    END p10
    PIN p11
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 13.405 51.555 13.475 ;
        END
    END p11
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 26.88 ;
      LAYER metal2 ;
        RECT  0 0 80.64 26.88 ;
      LAYER via1 ;
        RECT  0 0 80.64 26.88 ;
      LAYER metal1 ;
        RECT  0 0 80.64 26.88 ;
    END
END fake_macro_newblue1_o330113

MACRO fake_macro_newblue1_o330114
    CLASS BLOCK ;
    SIZE 80.64 BY 26.88 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 2.485 8.995 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 18.165 2.275 18.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.605 2.275 17.675 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 15.925 2.275 15.995 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.925 2.275 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 10.325 2.275 10.395 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 15.085 2.275 15.155 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 15.645 2.275 15.715 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 0.245 6.755 0.315 ;
        END
    END p9
    PIN p10
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.645 51.555 1.715 ;
        END
    END p10
    PIN p11
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 13.405 51.555 13.475 ;
        END
    END p11
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 26.88 ;
      LAYER metal2 ;
        RECT  0 0 80.64 26.88 ;
      LAYER via1 ;
        RECT  0 0 80.64 26.88 ;
      LAYER metal1 ;
        RECT  0 0 80.64 26.88 ;
    END
END fake_macro_newblue1_o330114

MACRO fake_macro_newblue1_o330115
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330115

MACRO fake_macro_newblue1_o330116
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330116

MACRO fake_macro_newblue1_o330117
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330117

MACRO fake_macro_newblue1_o330118
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330118

MACRO fake_macro_newblue1_o330119
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330119

MACRO fake_macro_newblue1_o330120
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330120

MACRO fake_macro_newblue1_o330121
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330121

MACRO fake_macro_newblue1_o330122
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330122

MACRO fake_macro_newblue1_o330123
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330123

MACRO fake_macro_newblue1_o330124
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330124

MACRO fake_macro_newblue1_o330125
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330125

MACRO fake_macro_newblue1_o330126
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330126

MACRO fake_macro_newblue1_o330127
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330127

MACRO fake_macro_newblue1_o330128
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330128

MACRO fake_macro_newblue1_o330129
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330129

MACRO fake_macro_newblue1_o330130
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330130

MACRO fake_macro_newblue1_o330131
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330131

MACRO fake_macro_newblue1_o330132
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330132

MACRO fake_macro_newblue1_o330133
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330133

MACRO fake_macro_newblue1_o330134
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330134

MACRO fake_macro_newblue1_o330135
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330135

MACRO fake_macro_newblue1_o330136
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330136

MACRO fake_macro_newblue1_o330137
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330137

MACRO fake_macro_newblue1_o330138
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330138

MACRO fake_macro_newblue1_o330139
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330139

MACRO fake_macro_newblue1_o330140
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330140

MACRO fake_macro_newblue1_o330141
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330141

MACRO fake_macro_newblue1_o330142
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330142

MACRO fake_macro_newblue1_o330143
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330143

MACRO fake_macro_newblue1_o330144
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330144

MACRO fake_macro_newblue1_o330145
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330145

MACRO fake_macro_newblue1_o330146
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330146

MACRO fake_macro_newblue1_o330147
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330147

MACRO fake_macro_newblue1_o330148
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330148

MACRO fake_macro_newblue1_o330149
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330149

MACRO fake_macro_newblue1_o330150
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330150

MACRO fake_macro_newblue1_o330151
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 73.605 0.035 73.675 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330151

MACRO fake_macro_newblue1_o330152
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330152

MACRO fake_macro_newblue1_o330153
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330153

MACRO fake_macro_newblue1_o330154
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330154

MACRO fake_macro_newblue1_o330155
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330155

MACRO fake_macro_newblue1_o330156
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330156

MACRO fake_macro_newblue1_o330157
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330157

MACRO fake_macro_newblue1_o330158
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330158

MACRO fake_macro_newblue1_o330159
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330159

MACRO fake_macro_newblue1_o330160
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330160

MACRO fake_macro_newblue1_o330161
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330161

MACRO fake_macro_newblue1_o330162
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330162

MACRO fake_macro_newblue1_o330163
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330163

MACRO fake_macro_newblue1_o330164
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330164

MACRO fake_macro_newblue1_o330165
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330165

MACRO fake_macro_newblue1_o330166
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330166

MACRO fake_macro_newblue1_o330167
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330167

MACRO fake_macro_newblue1_o330168
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330168

MACRO fake_macro_newblue1_o330169
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330169

MACRO fake_macro_newblue1_o330170
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330170

MACRO fake_macro_newblue1_o330171
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330171

MACRO fake_macro_newblue1_o330172
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330172

MACRO fake_macro_newblue1_o330173
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330173

MACRO fake_macro_newblue1_o330174
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330174

MACRO fake_macro_newblue1_o330175
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330175

MACRO fake_macro_newblue1_o330176
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330176

MACRO fake_macro_newblue1_o330177
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330177

MACRO fake_macro_newblue1_o330178
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330178

MACRO fake_macro_newblue1_o330179
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330179

MACRO fake_macro_newblue1_o330187
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330187

MACRO fake_macro_newblue1_o330188
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330188

MACRO fake_macro_newblue1_o330189
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330189

MACRO fake_macro_newblue1_o330190
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330190

MACRO fake_macro_newblue1_o330191
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330191

MACRO fake_macro_newblue1_o330192
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330192

MACRO fake_macro_newblue1_o330193
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330193

MACRO fake_macro_newblue1_o330194
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330194

MACRO fake_macro_newblue1_o330195
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330195

MACRO fake_macro_newblue1_o330196
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330196

MACRO fake_macro_newblue1_o330197
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330197

MACRO fake_macro_newblue1_o330198
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330198

MACRO fake_macro_newblue1_o330199
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330199

MACRO fake_macro_newblue1_o330200
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330200

MACRO fake_macro_newblue1_o330201
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330201

MACRO fake_macro_newblue1_o330202
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330202

MACRO fake_macro_newblue1_o330203
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330203

MACRO fake_macro_newblue1_o330204
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330204

MACRO fake_macro_newblue1_o330205
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330205

MACRO fake_macro_newblue1_o330206
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330206

MACRO fake_macro_newblue1_o330207
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330207

MACRO fake_macro_newblue1_o330208
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330208

MACRO fake_macro_newblue1_o330209
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330209

MACRO fake_macro_newblue1_o330210
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330210

MACRO fake_macro_newblue1_o330211
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330211

MACRO fake_macro_newblue1_o330212
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330212

MACRO fake_macro_newblue1_o330213
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 77.805 0.035 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 77.805 5.635 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.805 1.155 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 70.245 2.835 70.315 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330213

MACRO fake_macro_newblue1_o330214
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330214

MACRO fake_macro_newblue1_o330215
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330215

MACRO fake_macro_newblue1_o330216
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330216

MACRO fake_macro_newblue1_o330217
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330217

MACRO fake_macro_newblue1_o330218
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330218

MACRO fake_macro_newblue1_o330219
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330219

MACRO fake_macro_newblue1_o330220
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330220

MACRO fake_macro_newblue1_o330221
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330221

MACRO fake_macro_newblue1_o330222
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330222

MACRO fake_macro_newblue1_o330223
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330223

MACRO fake_macro_newblue1_o330224
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330224

MACRO fake_macro_newblue1_o330225
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330225

MACRO fake_macro_newblue1_o330226
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 12.845 77.875 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 7.245 77.875 7.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 11.725 77.875 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 10.045 77.875 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 13.125 73.395 13.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 10.045 70.035 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330226

MACRO fake_macro_newblue1_o330229
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330229

MACRO fake_macro_newblue1_o330230
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330230

MACRO fake_macro_newblue1_o330231
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330231

MACRO fake_macro_newblue1_o330232
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330232

MACRO fake_macro_newblue1_o330233
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330233

MACRO fake_macro_newblue1_o330234
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330234

MACRO fake_macro_newblue1_o330235
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330235

MACRO fake_macro_newblue1_o330236
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330236

MACRO fake_macro_newblue1_o330237
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330237

MACRO fake_macro_newblue1_o330238
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330238

MACRO fake_macro_newblue1_o330239
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330239

MACRO fake_macro_newblue1_o330240
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330240

MACRO fake_macro_newblue1_o330241
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330241

MACRO fake_macro_newblue1_o330242
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330242

MACRO fake_macro_newblue1_o330243
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330243

MACRO fake_macro_newblue1_o330244
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330244

MACRO fake_macro_newblue1_o330245
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330245

MACRO fake_macro_newblue1_o330246
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330246

MACRO fake_macro_newblue1_o330247
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330247

MACRO fake_macro_newblue1_o330248
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330248

MACRO fake_macro_newblue1_o330249
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330249

MACRO fake_macro_newblue1_o330250
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330250

MACRO fake_macro_newblue1_o330251
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330251

MACRO fake_macro_newblue1_o330252
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330252

MACRO fake_macro_newblue1_o330253
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330253

MACRO fake_macro_newblue1_o330254
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330254

MACRO fake_macro_newblue1_o330255
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330255

MACRO fake_macro_newblue1_o330256
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330256

MACRO fake_macro_newblue1_o330257
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330257

MACRO fake_macro_newblue1_o330258
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330258

MACRO fake_macro_newblue1_o330259
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330259

MACRO fake_macro_newblue1_o330260
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330260

MACRO fake_macro_newblue1_o330261
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330261

MACRO fake_macro_newblue1_o330262
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330262

MACRO fake_macro_newblue1_o330263
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330263

MACRO fake_macro_newblue1_o330264
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330264

MACRO fake_macro_newblue1_o330265
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330265

MACRO fake_macro_newblue1_o330266
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330266

MACRO fake_macro_newblue1_o330267
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330267

MACRO fake_macro_newblue1_o330268
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330268

MACRO fake_macro_newblue1_o330269
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330269

MACRO fake_macro_newblue1_o330270
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330270

MACRO fake_macro_newblue1_o330271
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330271

MACRO fake_macro_newblue1_o330272
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 2.485 12.355 2.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 2.485 5.075 2.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.485 9.555 2.555 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 2.485 10.675 2.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.685 12.355 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.045 9.555 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 51.765 12.915 51.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330272

MACRO fake_macro_newblue1_o330291
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330291

MACRO fake_macro_newblue1_o330292
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330292

MACRO fake_macro_newblue1_o330293
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330293

MACRO fake_macro_newblue1_o330294
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330294

MACRO fake_macro_newblue1_o330295
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330295

MACRO fake_macro_newblue1_o330296
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330296

MACRO fake_macro_newblue1_o330297
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330297

MACRO fake_macro_newblue1_o330298
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330298

MACRO fake_macro_newblue1_o330299
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330299

MACRO fake_macro_newblue1_o330300
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330300

MACRO fake_macro_newblue1_o330301
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330301

MACRO fake_macro_newblue1_o330302
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330302

MACRO fake_macro_newblue1_o330303
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330303

MACRO fake_macro_newblue1_o330304
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330304

MACRO fake_macro_newblue1_o330305
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330305

MACRO fake_macro_newblue1_o330306
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330306

MACRO fake_macro_newblue1_o330307
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330307

MACRO fake_macro_newblue1_o330308
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330308

MACRO fake_macro_newblue1_o330309
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330309

MACRO fake_macro_newblue1_o330310
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330310

MACRO fake_macro_newblue1_o330311
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330311

MACRO fake_macro_newblue1_o330312
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330312

MACRO fake_macro_newblue1_o330313
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330313

MACRO fake_macro_newblue1_o330314
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330314

MACRO fake_macro_newblue1_o330315
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330315

MACRO fake_macro_newblue1_o330316
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330316

MACRO fake_macro_newblue1_o330317
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330317

MACRO fake_macro_newblue1_o330318
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330318

MACRO fake_macro_newblue1_o330319
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330319

MACRO fake_macro_newblue1_o330320
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330320

MACRO fake_macro_newblue1_o330321
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330321

MACRO fake_macro_newblue1_o330322
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330322

MACRO fake_macro_newblue1_o330323
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330323

MACRO fake_macro_newblue1_o330324
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330324

MACRO fake_macro_newblue1_o330325
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330325

MACRO fake_macro_newblue1_o330326
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330326

MACRO fake_macro_newblue1_o330328
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330328

MACRO fake_macro_newblue1_o330329
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330329

MACRO fake_macro_newblue1_o330330
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330330

MACRO fake_macro_newblue1_o330331
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330331

MACRO fake_macro_newblue1_o330332
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330332

MACRO fake_macro_newblue1_o330333
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330333

MACRO fake_macro_newblue1_o330334
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330334

MACRO fake_macro_newblue1_o330335
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330335

MACRO fake_macro_newblue1_o330336
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330336

MACRO fake_macro_newblue1_o330337
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330337

MACRO fake_macro_newblue1_o330338
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330338

MACRO fake_macro_newblue1_o330339
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330339

MACRO fake_macro_newblue1_o330340
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330340

MACRO fake_macro_newblue1_o330341
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330341

MACRO fake_macro_newblue1_o330342
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330342

MACRO fake_macro_newblue1_o330343
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330343

MACRO fake_macro_newblue1_o330344
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330344

MACRO fake_macro_newblue1_o330345
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330345

MACRO fake_macro_newblue1_o330346
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330346

MACRO fake_macro_newblue1_o330347
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330347

MACRO fake_macro_newblue1_o330348
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330348

MACRO fake_macro_newblue1_o330349
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330349

MACRO fake_macro_newblue1_o330350
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330350

MACRO fake_macro_newblue1_o330351
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330351

MACRO fake_macro_newblue1_o330352
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330352

MACRO fake_macro_newblue1_o330353
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330353

MACRO fake_macro_newblue1_o330354
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330354

MACRO fake_macro_newblue1_o330355
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330355

MACRO fake_macro_newblue1_o330356
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330356

MACRO fake_macro_newblue1_o330357
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330357

MACRO fake_macro_newblue1_o330358
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330358

MACRO fake_macro_newblue1_o330359
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330359

MACRO fake_macro_newblue1_o330360
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330360

MACRO fake_macro_newblue1_o330361
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330361

MACRO fake_macro_newblue1_o330362
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330362

MACRO fake_macro_newblue1_o330363
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330363

MACRO fake_macro_newblue1_o330364
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330364

MACRO fake_macro_newblue1_o330365
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330365

MACRO fake_macro_newblue1_o330366
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330366

MACRO fake_macro_newblue1_o330367
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330367

MACRO fake_macro_newblue1_o330368
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330368

MACRO fake_macro_newblue1_o330369
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330369

MACRO fake_macro_newblue1_o330370
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330370

MACRO fake_macro_newblue1_o330371
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330371

MACRO fake_macro_newblue1_o330372
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 77.805 10.675 77.875 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330372

MACRO fake_macro_newblue1_o330373
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 10.885 2.275 10.955 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330373

MACRO fake_macro_newblue1_o330374
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 0.245 2.275 0.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.845 2.275 5.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.045 2.275 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 -0.035 6.755 0.035 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330374

MACRO fake_macro_newblue1_o330375
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330375

MACRO fake_macro_newblue1_o330376
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330376

MACRO fake_macro_newblue1_o330377
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330377

MACRO fake_macro_newblue1_o330378
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330378

MACRO fake_macro_newblue1_o330379
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330379

MACRO fake_macro_newblue1_o330380
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330380

MACRO fake_macro_newblue1_o330381
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330381

MACRO fake_macro_newblue1_o330382
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330382

MACRO fake_macro_newblue1_o330383
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330383

MACRO fake_macro_newblue1_o330384
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330384

MACRO fake_macro_newblue1_o330385
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 4.165 70.035 4.235 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330385

MACRO fake_macro_newblue1_o330386
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 8.085 77.875 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 0.805 77.875 0.875 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 9.205 77.875 9.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 2.765 73.395 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 13.125 28.595 13.195 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330386

MACRO fake_macro_newblue1_o330387
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330387

MACRO fake_macro_newblue1_o330388
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330388

MACRO fake_macro_newblue1_o330389
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330389

MACRO fake_macro_newblue1_o330390
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330390

MACRO fake_macro_newblue1_o330391
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330391

MACRO fake_macro_newblue1_o330392
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330392

MACRO fake_macro_newblue1_o330393
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330393

MACRO fake_macro_newblue1_o330394
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330394

MACRO fake_macro_newblue1_o330395
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330395

MACRO fake_macro_newblue1_o330396
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.005 2.275 12.075 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.845 2.275 12.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.005 2.275 5.075 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.285 2.275 12.355 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.885 2.275 3.955 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 10.325 6.755 10.395 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 8.925 10.115 8.995 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330396

MACRO fake_macro_newblue1_o330397
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330397

MACRO fake_macro_newblue1_o330398
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330398

MACRO fake_macro_newblue1_o330399
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330399

MACRO fake_macro_newblue1_o330400
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330400

MACRO fake_macro_newblue1_o330401
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330401

MACRO fake_macro_newblue1_o330402
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330402

MACRO fake_macro_newblue1_o330403
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330403

MACRO fake_macro_newblue1_o330404
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330404

MACRO fake_macro_newblue1_o330405
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330405

MACRO fake_macro_newblue1_o330406
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330406

MACRO fake_macro_newblue1_o330407
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330407

MACRO fake_macro_newblue1_o330408
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330408

MACRO fake_macro_newblue1_o330409
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330409

MACRO fake_macro_newblue1_o330410
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330410

MACRO fake_macro_newblue1_o330411
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330411

MACRO fake_macro_newblue1_o330412
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330412

MACRO fake_macro_newblue1_o330413
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330413

MACRO fake_macro_newblue1_o330414
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330414

MACRO fake_macro_newblue1_o330415
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330415

MACRO fake_macro_newblue1_o330416
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330416

MACRO fake_macro_newblue1_o330417
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330417

MACRO fake_macro_newblue1_o330418
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330418

MACRO fake_macro_newblue1_o330419
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330419

MACRO fake_macro_newblue1_o330420
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330420

MACRO fake_macro_newblue1_o330421
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330421

MACRO fake_macro_newblue1_o330422
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330422

MACRO fake_macro_newblue1_o330423
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330423

MACRO fake_macro_newblue1_o330424
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330424

MACRO fake_macro_newblue1_o330425
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330425

MACRO fake_macro_newblue1_o330426
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330426

MACRO fake_macro_newblue1_o330427
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330427

MACRO fake_macro_newblue1_o330428
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330428

MACRO fake_macro_newblue1_o330429
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.005 2.275 12.075 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.005 2.275 5.075 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.285 2.275 12.355 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.845 2.275 12.915 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.885 2.275 3.955 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 10.325 6.755 10.395 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 8.925 10.115 8.995 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330429

MACRO fake_macro_newblue1_o330430
    CLASS BLOCK ;
    SIZE 80.64 BY 13.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.005 2.275 12.075 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.845 2.275 12.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 5.005 2.275 5.075 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 12.285 2.275 12.355 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 3.885 2.275 3.955 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 10.325 6.755 10.395 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 8.925 10.115 8.995 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 -0.035 51.555 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal2 ;
        RECT  0 0 80.64 13.44 ;
      LAYER via1 ;
        RECT  0 0 80.64 13.44 ;
      LAYER metal1 ;
        RECT  0 0 80.64 13.44 ;
    END
END fake_macro_newblue1_o330430

MACRO fake_macro_newblue1_o330431
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330431

MACRO fake_macro_newblue1_o330432
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330432

MACRO fake_macro_newblue1_o330433
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330433

MACRO fake_macro_newblue1_o330434
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330434

MACRO fake_macro_newblue1_o330435
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330435

MACRO fake_macro_newblue1_o330436
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330436

MACRO fake_macro_newblue1_o330437
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330437

MACRO fake_macro_newblue1_o330438
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 70.245 8.995 70.315 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330438

MACRO fake_macro_newblue1_o330439
    CLASS BLOCK ;
    SIZE 13.44 BY 80.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 77.805 11.795 77.875 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 77.805 5.075 77.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 77.805 12.355 77.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 77.805 12.915 77.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 77.805 3.955 77.875 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 28.525 0.035 28.595 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal2 ;
        RECT  0 0 13.44 80.64 ;
      LAYER via1 ;
        RECT  0 0 13.44 80.64 ;
      LAYER metal1 ;
        RECT  0 0 13.44 80.64 ;
    END
END fake_macro_newblue1_o330439

MACRO fake_macro_newblue1_o330083
    CLASS BLOCK ;
    SIZE 838.04 BY 661.92 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  708.365 339.325 708.435 339.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 378.525 671.475 378.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 374.885 671.475 374.955 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 370.965 671.475 371.035 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 370.685 671.475 370.755 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 367.045 671.475 367.115 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 366.765 671.475 366.835 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 363.125 671.475 363.195 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 359.205 671.475 359.275 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 355.285 671.475 355.355 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 355.005 671.475 355.075 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 351.365 671.475 351.435 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 347.445 671.475 347.515 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 347.165 671.475 347.235 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 343.525 671.475 343.595 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 339.325 671.475 339.395 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 335.685 671.475 335.755 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 331.765 671.475 331.835 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 331.485 671.475 331.555 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 327.845 671.475 327.915 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 323.925 671.475 323.995 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 320.005 671.475 320.075 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  682.045 237.405 682.115 237.475 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  380.765 367.045 380.835 367.115 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 355.005 550.515 355.075 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 351.365 717.395 351.435 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 433.685 162.995 433.755 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 433.405 162.995 433.475 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 456.925 282.835 456.995 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 453.285 282.835 453.355 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 453.005 282.835 453.075 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 449.365 282.835 449.435 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 449.085 282.835 449.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 445.445 282.835 445.515 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 445.165 282.835 445.235 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 441.525 282.835 441.595 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 441.245 282.835 441.315 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 437.605 282.835 437.675 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 437.325 282.835 437.395 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 433.685 282.835 433.755 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 433.405 282.835 433.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 429.765 282.835 429.835 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 429.485 282.835 429.555 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 425.845 282.835 425.915 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 425.565 282.835 425.635 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 421.925 282.835 421.995 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 421.645 282.835 421.715 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 418.005 282.835 418.075 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 417.725 282.835 417.795 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 414.085 282.835 414.155 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 413.805 282.835 413.875 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 410.165 282.835 410.235 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 409.885 282.835 409.955 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 406.245 282.835 406.315 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 405.965 282.835 406.035 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 402.325 282.835 402.395 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 402.045 282.835 402.115 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 398.405 282.835 398.475 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 398.125 282.835 398.195 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  282.765 394.485 282.835 394.555 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 456.925 248.115 456.995 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 453.285 248.115 453.355 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 453.005 248.115 453.075 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 449.365 248.115 449.435 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 449.085 248.115 449.155 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 445.445 248.115 445.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 445.165 248.115 445.235 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 441.525 248.115 441.595 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 441.245 248.115 441.315 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 437.605 248.115 437.675 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 437.325 248.115 437.395 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 433.685 248.115 433.755 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 433.405 248.115 433.475 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 429.765 248.115 429.835 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 429.485 248.115 429.555 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 425.845 248.115 425.915 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 425.565 248.115 425.635 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 421.925 248.115 421.995 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 421.645 248.115 421.715 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 418.005 248.115 418.075 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 417.725 248.115 417.795 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 414.085 248.115 414.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 413.805 248.115 413.875 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 410.165 248.115 410.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 409.885 248.115 409.955 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 406.245 248.115 406.315 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 405.965 248.115 406.035 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 402.325 248.115 402.395 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 402.045 248.115 402.115 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 398.405 248.115 398.475 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 398.125 248.115 398.195 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 394.485 248.115 394.555 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 429.765 162.995 429.835 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 300.125 251.475 300.195 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 296.485 251.475 296.555 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 296.205 251.475 296.275 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 292.565 251.475 292.635 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 292.285 251.475 292.355 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 288.645 251.475 288.715 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 288.365 251.475 288.435 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 284.725 251.475 284.795 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 284.445 251.475 284.515 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 280.805 251.475 280.875 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 280.525 251.475 280.595 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 276.885 251.475 276.955 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 276.605 251.475 276.675 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 272.965 251.475 273.035 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 272.685 251.475 272.755 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 269.045 251.475 269.115 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 268.765 251.475 268.835 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 265.125 251.475 265.195 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 264.845 251.475 264.915 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 261.205 251.475 261.275 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 260.925 251.475 260.995 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 257.285 251.475 257.355 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 257.005 251.475 257.075 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 253.365 251.475 253.435 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 253.085 251.475 253.155 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 249.445 251.475 249.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 249.165 251.475 249.235 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 245.525 251.475 245.595 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 245.245 251.475 245.315 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 241.605 251.475 241.675 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 241.325 251.475 241.395 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  251.405 237.685 251.475 237.755 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  224.525 319.725 224.595 319.795 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  224.525 320.005 224.595 320.075 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  259.805 315.805 259.875 315.875 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 366.765 717.395 366.835 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 363.125 717.395 363.195 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  380.765 366.765 380.835 366.835 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 351.085 550.515 351.155 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 347.445 550.515 347.515 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 359.205 550.515 359.275 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 323.645 550.515 323.715 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 323.925 550.515 323.995 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  492.205 300.125 492.275 300.195 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 296.485 493.395 296.555 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  492.765 296.205 492.835 296.275 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  489.405 292.565 489.475 292.635 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 292.285 493.395 292.355 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 288.645 493.395 288.715 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  488.285 288.365 488.355 288.435 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 284.725 493.395 284.795 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 284.445 493.395 284.515 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 280.805 493.395 280.875 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  487.725 280.525 487.795 280.595 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 276.885 486.115 276.955 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 276.605 493.395 276.675 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 272.965 493.395 273.035 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  492.205 272.685 492.275 272.755 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 269.325 486.115 269.395 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 268.765 486.115 268.835 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 265.125 486.115 265.195 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 264.845 486.115 264.915 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  492.205 261.205 492.275 261.275 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 260.925 486.115 260.995 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  493.325 257.285 493.395 257.355 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 257.285 486.115 257.355 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 253.645 486.115 253.715 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 252.525 486.115 252.595 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  492.205 249.445 492.275 249.515 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 249.165 486.115 249.235 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 245.805 486.115 245.875 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 245.245 486.115 245.315 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 241.325 486.115 241.395 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  492.205 241.325 492.275 241.395 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  486.045 237.685 486.115 237.755 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  544.285 351.365 544.355 351.435 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 378.805 550.515 378.875 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  535.885 374.325 535.955 374.395 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  546.525 370.965 546.595 371.035 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  544.285 370.685 544.355 370.755 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  568.925 296.485 568.995 296.555 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  568.925 324.205 568.995 324.275 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  568.925 296.205 568.995 296.275 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  568.925 295.925 568.995 295.995 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  503.405 339.605 503.475 339.675 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  505.085 339.605 505.155 339.675 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 367.045 550.515 367.115 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 327.565 550.515 327.635 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 327.845 550.515 327.915 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 366.765 550.515 366.835 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 339.325 550.515 339.395 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 331.485 550.515 331.555 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 331.765 550.515 331.835 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 362.845 550.515 362.915 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 350.805 550.515 350.875 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 347.165 550.515 347.235 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  551.005 324.205 551.075 324.275 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 358.925 550.515 358.995 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  515.165 331.485 515.235 331.555 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  515.165 327.565 515.235 327.635 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  515.165 331.765 515.235 331.835 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  515.165 327.845 515.235 327.915 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  515.165 335.405 515.235 335.475 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 343.525 550.515 343.595 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 355.285 550.515 355.355 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 335.405 550.515 335.475 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 335.685 550.515 335.755 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  550.445 374.885 550.515 374.955 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  551.005 332.045 551.075 332.115 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 488.285 117.075 488.355 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 437.325 162.995 437.395 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  187.005 300.405 187.075 300.475 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 182.525 159.635 182.595 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  287.805 237.685 287.875 237.755 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  313.005 367.045 313.075 367.115 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  287.245 449.365 287.315 449.435 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  273.245 457.205 273.315 457.275 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  367.885 496.125 367.955 496.195 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  350.525 453.005 350.595 453.075 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 174.965 330.435 175.035 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  387.485 123.725 387.555 123.795 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  387.485 190.365 387.555 190.435 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  387.485 229.845 387.555 229.915 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  385.805 433.685 385.875 433.755 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  476.525 449.365 476.595 449.435 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 382.445 671.475 382.515 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 378.805 671.475 378.875 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 374.605 671.475 374.675 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 362.845 671.475 362.915 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 358.925 671.475 358.995 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 351.085 671.475 351.155 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 343.245 671.475 343.315 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 339.605 671.475 339.675 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 335.405 671.475 335.475 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 327.565 671.475 327.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 323.645 671.475 323.715 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 335.685 717.395 335.755 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 358.925 330.435 358.995 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 351.085 717.395 351.155 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 366.765 330.435 366.835 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 421.645 162.995 421.715 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 233.765 133.315 233.835 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 437.605 162.995 437.675 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 425.565 162.995 425.635 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 398.125 162.995 398.195 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 445.445 162.995 445.515 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 480.445 280.035 480.515 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 508.165 280.035 508.235 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 480.725 280.035 480.795 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  280.525 481.005 280.595 481.075 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 484.365 280.035 484.435 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  280.525 484.645 280.595 484.715 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 484.645 280.035 484.715 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  280.525 484.925 280.595 484.995 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 488.285 280.035 488.355 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  280.525 488.565 280.595 488.635 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 488.565 280.035 488.635 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  280.525 488.845 280.595 488.915 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 492.205 280.035 492.275 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  280.525 492.485 280.595 492.555 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  279.965 492.485 280.035 492.555 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  280.525 492.765 280.595 492.835 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 480.445 315.315 480.515 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 508.165 315.315 508.235 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 480.725 315.315 480.795 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.805 481.005 315.875 481.075 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 484.365 315.315 484.435 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.805 484.645 315.875 484.715 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 484.645 315.315 484.715 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.805 484.925 315.875 484.995 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 488.285 315.315 488.355 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.805 488.565 315.875 488.635 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 488.565 315.315 488.635 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.805 488.845 315.875 488.915 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 492.205 315.315 492.275 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.805 492.485 315.875 492.555 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.245 492.485 315.315 492.555 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  315.805 492.765 315.875 492.835 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 480.445 402.675 480.515 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 508.165 402.675 508.235 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 480.725 402.675 480.795 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  403.165 481.005 403.235 481.075 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 484.365 402.675 484.435 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  403.165 484.645 403.235 484.715 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 484.645 402.675 484.715 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  403.165 484.925 403.235 484.995 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 488.285 402.675 488.355 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  403.165 488.565 403.235 488.635 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 488.565 402.675 488.635 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  403.165 488.845 403.235 488.915 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 492.205 402.675 492.275 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  403.165 492.485 403.235 492.555 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  402.605 492.485 402.675 492.555 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  403.165 492.765 403.235 492.835 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 480.445 437.955 480.515 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 508.165 437.955 508.235 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 480.725 437.955 480.795 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  438.445 481.005 438.515 481.075 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 484.365 437.955 484.435 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  438.445 484.645 438.515 484.715 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 484.645 437.955 484.715 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  438.445 484.925 438.515 484.995 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 488.285 437.955 488.355 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  438.445 488.565 438.515 488.635 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 488.565 437.955 488.635 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  438.445 488.845 438.515 488.915 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 492.205 437.955 492.275 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  438.445 492.485 438.515 492.555 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  437.885 492.485 437.955 492.555 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  438.445 492.765 438.515 492.835 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  142.205 159.285 142.275 159.355 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  142.205 187.005 142.275 187.075 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.925 159.285 106.995 159.355 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 159.285 71.715 159.355 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 187.005 71.715 187.075 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 159.285 36.435 159.355 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 159.285 1.715 159.355 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 187.005 1.715 187.075 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  142.205 159.005 142.275 159.075 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.925 159.005 106.995 159.075 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.925 186.725 106.995 186.795 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 159.005 71.715 159.075 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 158.725 71.715 158.795 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 159.005 36.435 159.075 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 186.725 36.435 186.795 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 159.005 1.715 159.075 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.085 229.565 169.155 229.635 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.085 257.285 169.155 257.355 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.085 229.845 169.155 229.915 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.645 230.125 169.715 230.195 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.085 233.485 169.155 233.555 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.645 233.765 169.715 233.835 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.085 233.765 169.155 233.835 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.645 234.045 169.715 234.115 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 398.405 162.995 398.475 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  248.045 394.205 248.115 394.275 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  224.525 323.645 224.595 323.715 ;
        END
    END p329
    PIN p330
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 441.245 162.995 441.315 ;
        END
    END p330
    PIN p331
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 362.845 330.435 362.915 ;
        END
    END p331
    PIN p332
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  353.885 375.445 353.955 375.515 ;
        END
    END p332
    PIN p333
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  380.765 358.925 380.835 358.995 ;
        END
    END p333
    PIN p334
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  380.765 363.125 380.835 363.195 ;
        END
    END p334
    PIN p335
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  380.765 362.845 380.835 362.915 ;
        END
    END p335
    PIN p336
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  380.765 359.205 380.835 359.275 ;
        END
    END p336
    PIN p337
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 362.845 717.395 362.915 ;
        END
    END p337
    PIN p338
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 367.045 717.395 367.115 ;
        END
    END p338
    PIN p339
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 320.005 619.955 320.075 ;
        END
    END p339
    PIN p340
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 323.645 619.955 323.715 ;
        END
    END p340
    PIN p341
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 323.925 619.955 323.995 ;
        END
    END p341
    PIN p342
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 327.565 619.955 327.635 ;
        END
    END p342
    PIN p343
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 327.845 619.955 327.915 ;
        END
    END p343
    PIN p344
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 331.485 619.955 331.555 ;
        END
    END p344
    PIN p345
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 331.765 619.955 331.835 ;
        END
    END p345
    PIN p346
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 335.405 619.955 335.475 ;
        END
    END p346
    PIN p347
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 335.685 619.955 335.755 ;
        END
    END p347
    PIN p348
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 339.325 619.955 339.395 ;
        END
    END p348
    PIN p349
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 339.605 619.955 339.675 ;
        END
    END p349
    PIN p350
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 343.245 619.955 343.315 ;
        END
    END p350
    PIN p351
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 343.525 619.955 343.595 ;
        END
    END p351
    PIN p352
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 347.165 619.955 347.235 ;
        END
    END p352
    PIN p353
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 347.445 619.955 347.515 ;
        END
    END p353
    PIN p354
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 351.085 619.955 351.155 ;
        END
    END p354
    PIN p355
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 351.365 619.955 351.435 ;
        END
    END p355
    PIN p356
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 355.005 619.955 355.075 ;
        END
    END p356
    PIN p357
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 355.285 619.955 355.355 ;
        END
    END p357
    PIN p358
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 358.925 619.955 358.995 ;
        END
    END p358
    PIN p359
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 359.205 619.955 359.275 ;
        END
    END p359
    PIN p360
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 362.845 619.955 362.915 ;
        END
    END p360
    PIN p361
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 363.125 619.955 363.195 ;
        END
    END p361
    PIN p362
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 366.765 619.955 366.835 ;
        END
    END p362
    PIN p363
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 367.045 619.955 367.115 ;
        END
    END p363
    PIN p364
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 370.685 619.955 370.755 ;
        END
    END p364
    PIN p365
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 370.965 619.955 371.035 ;
        END
    END p365
    PIN p366
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 374.605 619.955 374.675 ;
        END
    END p366
    PIN p367
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 374.885 619.955 374.955 ;
        END
    END p367
    PIN p368
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 378.525 619.955 378.595 ;
        END
    END p368
    PIN p369
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 378.805 619.955 378.875 ;
        END
    END p369
    PIN p370
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 382.445 619.955 382.515 ;
        END
    END p370
    PIN p371
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 379.085 717.395 379.155 ;
        END
    END p371
    PIN p372
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  707.245 355.285 707.315 355.355 ;
        END
    END p372
    PIN p373
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 355.005 717.395 355.075 ;
        END
    END p373
    PIN p374
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  716.765 327.845 716.835 327.915 ;
        END
    END p374
    PIN p375
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 331.485 717.395 331.555 ;
        END
    END p375
    PIN p376
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 331.765 717.395 331.835 ;
        END
    END p376
    PIN p377
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 359.205 330.435 359.275 ;
        END
    END p377
    PIN p378
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 386.645 330.435 386.715 ;
        END
    END p378
    PIN p379
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  224.525 331.485 224.595 331.555 ;
        END
    END p379
    PIN p380
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  224.525 327.845 224.595 327.915 ;
        END
    END p380
    PIN p381
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 363.125 330.435 363.195 ;
        END
    END p381
    PIN p382
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  220.605 374.885 220.675 374.955 ;
        END
    END p382
    PIN p383
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  202.685 374.885 202.755 374.955 ;
        END
    END p383
    PIN p384
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  435.085 194.565 435.155 194.635 ;
        END
    END p384
    PIN p385
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 328.405 702.275 328.475 ;
        END
    END p385
    PIN p386
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  435.085 194.285 435.155 194.355 ;
        END
    END p386
    PIN p387
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  247.485 178.885 247.555 178.955 ;
        END
    END p387
    PIN p388
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  246.925 178.885 246.995 178.955 ;
        END
    END p388
    PIN p389
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  212.205 178.885 212.275 178.955 ;
        END
    END p389
    PIN p390
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  212.205 206.605 212.275 206.675 ;
        END
    END p390
    PIN p391
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  176.925 178.885 176.995 178.955 ;
        END
    END p391
    PIN p392
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  176.925 206.605 176.995 206.675 ;
        END
    END p392
    PIN p393
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  142.205 178.885 142.275 178.955 ;
        END
    END p393
    PIN p394
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  142.765 179.165 142.835 179.235 ;
        END
    END p394
    PIN p395
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.925 178.885 106.995 178.955 ;
        END
    END p395
    PIN p396
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  107.485 179.165 107.555 179.235 ;
        END
    END p396
    PIN p397
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 178.885 71.715 178.955 ;
        END
    END p397
    PIN p398
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.205 179.165 72.275 179.235 ;
        END
    END p398
    PIN p399
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 178.885 36.435 178.955 ;
        END
    END p399
    PIN p400
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 179.165 36.995 179.235 ;
        END
    END p400
    PIN p401
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 178.885 1.715 178.955 ;
        END
    END p401
    PIN p402
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 179.165 2.275 179.235 ;
        END
    END p402
    PIN p403
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  554.925 178.885 554.995 178.955 ;
        END
    END p403
    PIN p404
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  554.925 206.605 554.995 206.675 ;
        END
    END p404
    PIN p405
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  590.205 178.885 590.275 178.955 ;
        END
    END p405
    PIN p406
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  590.205 206.605 590.275 206.675 ;
        END
    END p406
    PIN p407
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  625.485 178.885 625.555 178.955 ;
        END
    END p407
    PIN p408
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  625.485 206.605 625.555 206.675 ;
        END
    END p408
    PIN p409
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  660.765 178.885 660.835 178.955 ;
        END
    END p409
    PIN p410
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  660.765 206.605 660.835 206.675 ;
        END
    END p410
    PIN p411
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  695.485 178.885 695.555 178.955 ;
        END
    END p411
    PIN p412
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  695.485 206.605 695.555 206.675 ;
        END
    END p412
    PIN p413
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  730.765 178.885 730.835 178.955 ;
        END
    END p413
    PIN p414
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  730.765 206.605 730.835 206.675 ;
        END
    END p414
    PIN p415
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  766.045 178.885 766.115 178.955 ;
        END
    END p415
    PIN p416
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  766.045 206.605 766.115 206.675 ;
        END
    END p416
    PIN p417
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  801.325 178.885 801.395 178.955 ;
        END
    END p417
    PIN p418
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  801.325 206.605 801.395 206.675 ;
        END
    END p418
    PIN p419
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  247.485 178.605 247.555 178.675 ;
        END
    END p419
    PIN p420
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  246.925 178.605 246.995 178.675 ;
        END
    END p420
    PIN p421
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  212.205 178.605 212.275 178.675 ;
        END
    END p421
    PIN p422
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 178.325 208.355 178.395 ;
        END
    END p422
    PIN p423
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  176.925 178.605 176.995 178.675 ;
        END
    END p423
    PIN p424
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  176.925 178.325 176.995 178.395 ;
        END
    END p424
    PIN p425
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  142.205 178.605 142.275 178.675 ;
        END
    END p425
    PIN p426
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  139.405 178.325 139.475 178.395 ;
        END
    END p426
    PIN p427
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.925 178.605 106.995 178.675 ;
        END
    END p427
    PIN p428
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  107.485 178.885 107.555 178.955 ;
        END
    END p428
    PIN p429
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 178.605 71.715 178.675 ;
        END
    END p429
    PIN p430
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.205 178.885 72.275 178.955 ;
        END
    END p430
    PIN p431
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 178.605 36.435 178.675 ;
        END
    END p431
    PIN p432
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 178.885 36.995 178.955 ;
        END
    END p432
    PIN p433
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 178.605 1.715 178.675 ;
        END
    END p433
    PIN p434
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 178.885 2.275 178.955 ;
        END
    END p434
    PIN p435
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  554.925 178.605 554.995 178.675 ;
        END
    END p435
    PIN p436
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  554.925 178.325 554.995 178.395 ;
        END
    END p436
    PIN p437
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  590.205 178.605 590.275 178.675 ;
        END
    END p437
    PIN p438
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  590.205 178.325 590.275 178.395 ;
        END
    END p438
    PIN p439
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  625.485 178.605 625.555 178.675 ;
        END
    END p439
    PIN p440
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  625.485 178.325 625.555 178.395 ;
        END
    END p440
    PIN p441
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  660.765 178.605 660.835 178.675 ;
        END
    END p441
    PIN p442
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  660.765 178.325 660.835 178.395 ;
        END
    END p442
    PIN p443
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  695.485 178.605 695.555 178.675 ;
        END
    END p443
    PIN p444
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  695.485 178.325 695.555 178.395 ;
        END
    END p444
    PIN p445
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  730.765 178.605 730.835 178.675 ;
        END
    END p445
    PIN p446
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  730.765 178.325 730.835 178.395 ;
        END
    END p446
    PIN p447
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  766.045 178.605 766.115 178.675 ;
        END
    END p447
    PIN p448
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  766.045 178.325 766.115 178.395 ;
        END
    END p448
    PIN p449
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  801.325 178.605 801.395 178.675 ;
        END
    END p449
    PIN p450
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  801.325 178.325 801.395 178.395 ;
        END
    END p450
    PIN p451
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  435.085 178.605 435.155 178.675 ;
        END
    END p451
    PIN p452
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  435.085 206.325 435.155 206.395 ;
        END
    END p452
    PIN p453
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  435.085 178.885 435.155 178.955 ;
        END
    END p453
    PIN p454
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  435.645 194.845 435.715 194.915 ;
        END
    END p454
    PIN p455
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  435.645 194.565 435.715 194.635 ;
        END
    END p455
    PIN p456
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 441.525 162.995 441.595 ;
        END
    END p456
    PIN p457
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 445.165 162.995 445.235 ;
        END
    END p457
    PIN p458
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 449.085 162.995 449.155 ;
        END
    END p458
    PIN p459
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 449.365 162.995 449.435 ;
        END
    END p459
    PIN p460
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 453.005 162.995 453.075 ;
        END
    END p460
    PIN p461
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 350.805 717.395 350.875 ;
        END
    END p461
    PIN p462
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.885 332.045 717.955 332.115 ;
        END
    END p462
    PIN p463
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 335.405 717.395 335.475 ;
        END
    END p463
    PIN p464
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  711.165 362.845 711.235 362.915 ;
        END
    END p464
    PIN p465
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  701.085 339.885 701.155 339.955 ;
        END
    END p465
    PIN p466
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 320.005 459.235 320.075 ;
        END
    END p466
    PIN p467
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 323.645 459.235 323.715 ;
        END
    END p467
    PIN p468
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 323.925 459.235 323.995 ;
        END
    END p468
    PIN p469
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 327.565 459.235 327.635 ;
        END
    END p469
    PIN p470
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 327.845 459.235 327.915 ;
        END
    END p470
    PIN p471
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 331.485 459.235 331.555 ;
        END
    END p471
    PIN p472
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 331.765 459.235 331.835 ;
        END
    END p472
    PIN p473
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 335.405 459.235 335.475 ;
        END
    END p473
    PIN p474
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 335.685 459.235 335.755 ;
        END
    END p474
    PIN p475
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  459.165 339.325 459.235 339.395 ;
        END
    END p475
    PIN p476
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  701.645 394.485 701.715 394.555 ;
        END
    END p476
    PIN p477
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  713.965 398.125 714.035 398.195 ;
        END
    END p477
    PIN p478
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  701.645 398.685 701.715 398.755 ;
        END
    END p478
    PIN p479
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  715.645 402.045 715.715 402.115 ;
        END
    END p479
    PIN p480
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  716.765 402.325 716.835 402.395 ;
        END
    END p480
    PIN p481
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 405.965 717.395 406.035 ;
        END
    END p481
    PIN p482
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 406.245 717.395 406.315 ;
        END
    END p482
    PIN p483
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  701.085 409.885 701.155 409.955 ;
        END
    END p483
    PIN p484
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 410.445 702.275 410.515 ;
        END
    END p484
    PIN p485
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  701.085 413.525 701.155 413.595 ;
        END
    END p485
    PIN p486
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 414.085 702.275 414.155 ;
        END
    END p486
    PIN p487
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  716.765 417.725 716.835 417.795 ;
        END
    END p487
    PIN p488
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 418.285 702.275 418.355 ;
        END
    END p488
    PIN p489
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 421.645 702.275 421.715 ;
        END
    END p489
    PIN p490
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  716.765 421.925 716.835 421.995 ;
        END
    END p490
    PIN p491
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  701.645 425.565 701.715 425.635 ;
        END
    END p491
    PIN p492
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  713.965 425.845 714.035 425.915 ;
        END
    END p492
    PIN p493
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 429.205 702.275 429.275 ;
        END
    END p493
    PIN p494
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  713.965 429.765 714.035 429.835 ;
        END
    END p494
    PIN p495
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 433.405 717.395 433.475 ;
        END
    END p495
    PIN p496
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  716.765 433.685 716.835 433.755 ;
        END
    END p496
    PIN p497
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 437.325 702.275 437.395 ;
        END
    END p497
    PIN p498
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 437.605 702.275 437.675 ;
        END
    END p498
    PIN p499
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 441.245 717.395 441.315 ;
        END
    END p499
    PIN p500
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 441.525 717.395 441.595 ;
        END
    END p500
    PIN p501
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 445.165 702.275 445.235 ;
        END
    END p501
    PIN p502
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 445.445 717.395 445.515 ;
        END
    END p502
    PIN p503
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 448.805 702.275 448.875 ;
        END
    END p503
    PIN p504
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 449.925 702.275 449.995 ;
        END
    END p504
    PIN p505
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 452.445 702.275 452.515 ;
        END
    END p505
    PIN p506
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 453.005 702.275 453.075 ;
        END
    END p506
    PIN p507
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 457.205 702.275 457.275 ;
        END
    END p507
    PIN p508
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  712.845 366.765 712.915 366.835 ;
        END
    END p508
    PIN p509
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  702.205 367.325 702.275 367.395 ;
        END
    END p509
    PIN p510
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 347.165 717.395 347.235 ;
        END
    END p510
    PIN p511
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 347.445 717.395 347.515 ;
        END
    END p511
    PIN p512
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  169.085 300.125 169.155 300.195 ;
        END
    END p512
    PIN p513
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 111.685 330.435 111.755 ;
        END
    END p513
    PIN p514
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  430.605 398.125 430.675 398.195 ;
        END
    END p514
    PIN p515
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  515.165 343.245 515.235 343.315 ;
        END
    END p515
    PIN p516
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  510.685 155.085 510.755 155.155 ;
        END
    END p516
    PIN p517
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  568.925 260.925 568.995 260.995 ;
        END
    END p517
    PIN p518
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  618.205 319.725 618.275 319.795 ;
        END
    END p518
    PIN p519
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 402.325 619.955 402.395 ;
        END
    END p519
    PIN p520
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  619.885 441.525 619.955 441.595 ;
        END
    END p520
    PIN p521
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 449.085 671.475 449.155 ;
        END
    END p521
    PIN p522
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  671.405 402.325 671.475 402.395 ;
        END
    END p522
    PIN p523
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  682.045 251.125 682.115 251.195 ;
        END
    END p523
    PIN p524
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  695.485 155.085 695.555 155.155 ;
        END
    END p524
    PIN p525
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 421.645 26.355 421.715 ;
        END
    END p525
    PIN p526
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 253.365 52.675 253.435 ;
        END
    END p526
    PIN p527
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 237.405 133.315 237.475 ;
        END
    END p527
    PIN p528
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 347.445 117.075 347.515 ;
        END
    END p528
    PIN p529
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 233.765 330.435 233.835 ;
        END
    END p529
    PIN p530
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 237.685 204.435 237.755 ;
        END
    END p530
    PIN p531
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 241.325 204.435 241.395 ;
        END
    END p531
    PIN p532
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 241.605 204.435 241.675 ;
        END
    END p532
    PIN p533
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 245.245 204.435 245.315 ;
        END
    END p533
    PIN p534
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 245.525 204.435 245.595 ;
        END
    END p534
    PIN p535
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 249.165 204.435 249.235 ;
        END
    END p535
    PIN p536
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 249.445 204.435 249.515 ;
        END
    END p536
    PIN p537
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 253.085 204.435 253.155 ;
        END
    END p537
    PIN p538
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 253.365 204.435 253.435 ;
        END
    END p538
    PIN p539
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 257.005 204.435 257.075 ;
        END
    END p539
    PIN p540
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 257.285 204.435 257.355 ;
        END
    END p540
    PIN p541
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 260.925 204.435 260.995 ;
        END
    END p541
    PIN p542
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 261.205 204.435 261.275 ;
        END
    END p542
    PIN p543
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 264.845 204.435 264.915 ;
        END
    END p543
    PIN p544
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 265.125 204.435 265.195 ;
        END
    END p544
    PIN p545
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 268.765 204.435 268.835 ;
        END
    END p545
    PIN p546
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 269.045 204.435 269.115 ;
        END
    END p546
    PIN p547
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 272.685 204.435 272.755 ;
        END
    END p547
    PIN p548
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 272.965 204.435 273.035 ;
        END
    END p548
    PIN p549
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 276.605 204.435 276.675 ;
        END
    END p549
    PIN p550
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 276.885 204.435 276.955 ;
        END
    END p550
    PIN p551
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 280.525 204.435 280.595 ;
        END
    END p551
    PIN p552
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 280.805 204.435 280.875 ;
        END
    END p552
    PIN p553
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 284.445 204.435 284.515 ;
        END
    END p553
    PIN p554
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 284.725 204.435 284.795 ;
        END
    END p554
    PIN p555
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 288.365 204.435 288.435 ;
        END
    END p555
    PIN p556
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 288.645 204.435 288.715 ;
        END
    END p556
    PIN p557
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 292.285 204.435 292.355 ;
        END
    END p557
    PIN p558
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 292.565 204.435 292.635 ;
        END
    END p558
    PIN p559
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 296.205 204.435 296.275 ;
        END
    END p559
    PIN p560
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 296.485 204.435 296.555 ;
        END
    END p560
    PIN p561
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  204.365 300.125 204.435 300.195 ;
        END
    END p561
    PIN p562
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 229.565 133.315 229.635 ;
        END
    END p562
    PIN p563
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 261.485 330.435 261.555 ;
        END
    END p563
    PIN p564
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  330.365 233.485 330.435 233.555 ;
        END
    END p564
    PIN p565
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 233.485 133.315 233.555 ;
        END
    END p565
    PIN p566
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  247.485 159.285 247.555 159.355 ;
        END
    END p566
    PIN p567
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  247.485 187.005 247.555 187.075 ;
        END
    END p567
    PIN p568
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  212.205 159.285 212.275 159.355 ;
        END
    END p568
    PIN p569
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  212.205 178.325 212.275 178.395 ;
        END
    END p569
    PIN p570
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  176.925 159.285 176.995 159.355 ;
        END
    END p570
    PIN p571
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  177.485 159.565 177.555 159.635 ;
        END
    END p571
    PIN p572
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  107.485 159.565 107.555 159.635 ;
        END
    END p572
    PIN p573
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 159.565 36.995 159.635 ;
        END
    END p573
    PIN p574
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  554.925 159.285 554.995 159.355 ;
        END
    END p574
    PIN p575
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  555.485 159.565 555.555 159.635 ;
        END
    END p575
    PIN p576
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  590.205 159.285 590.275 159.355 ;
        END
    END p576
    PIN p577
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  590.765 159.565 590.835 159.635 ;
        END
    END p577
    PIN p578
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  625.485 159.285 625.555 159.355 ;
        END
    END p578
    PIN p579
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  626.045 159.565 626.115 159.635 ;
        END
    END p579
    PIN p580
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  660.765 159.285 660.835 159.355 ;
        END
    END p580
    PIN p581
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  661.325 159.565 661.395 159.635 ;
        END
    END p581
    PIN p582
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  695.485 159.285 695.555 159.355 ;
        END
    END p582
    PIN p583
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  696.045 159.565 696.115 159.635 ;
        END
    END p583
    PIN p584
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  730.765 159.285 730.835 159.355 ;
        END
    END p584
    PIN p585
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  731.325 159.565 731.395 159.635 ;
        END
    END p585
    PIN p586
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  766.045 159.285 766.115 159.355 ;
        END
    END p586
    PIN p587
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  766.605 159.565 766.675 159.635 ;
        END
    END p587
    PIN p588
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  801.325 159.285 801.395 159.355 ;
        END
    END p588
    PIN p589
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  801.885 159.565 801.955 159.635 ;
        END
    END p589
    PIN p590
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  247.485 159.005 247.555 159.075 ;
        END
    END p590
    PIN p591
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  247.485 158.725 247.555 158.795 ;
        END
    END p591
    PIN p592
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  212.205 159.005 212.275 159.075 ;
        END
    END p592
    PIN p593
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  212.205 158.725 212.275 158.795 ;
        END
    END p593
    PIN p594
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  176.925 159.005 176.995 159.075 ;
        END
    END p594
    PIN p595
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  177.485 159.285 177.555 159.355 ;
        END
    END p595
    PIN p596
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  142.205 158.725 142.275 158.795 ;
        END
    END p596
    PIN p597
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 159.285 2.275 159.355 ;
        END
    END p597
    PIN p598
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  554.925 159.005 554.995 159.075 ;
        END
    END p598
    PIN p599
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  555.485 159.285 555.555 159.355 ;
        END
    END p599
    PIN p600
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  590.205 159.005 590.275 159.075 ;
        END
    END p600
    PIN p601
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  590.765 159.285 590.835 159.355 ;
        END
    END p601
    PIN p602
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  625.485 159.005 625.555 159.075 ;
        END
    END p602
    PIN p603
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  626.045 159.285 626.115 159.355 ;
        END
    END p603
    PIN p604
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  660.765 159.005 660.835 159.075 ;
        END
    END p604
    PIN p605
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  661.325 159.285 661.395 159.355 ;
        END
    END p605
    PIN p606
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  695.485 159.005 695.555 159.075 ;
        END
    END p606
    PIN p607
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  696.045 159.285 696.115 159.355 ;
        END
    END p607
    PIN p608
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  730.765 159.005 730.835 159.075 ;
        END
    END p608
    PIN p609
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  731.325 159.285 731.395 159.355 ;
        END
    END p609
    PIN p610
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  766.045 159.005 766.115 159.075 ;
        END
    END p610
    PIN p611
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  766.605 159.285 766.675 159.355 ;
        END
    END p611
    PIN p612
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  801.325 159.005 801.395 159.075 ;
        END
    END p612
    PIN p613
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  801.885 159.285 801.955 159.355 ;
        END
    END p613
    PIN p614
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 394.485 208.355 394.555 ;
        END
    END p614
    PIN p615
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 398.125 208.355 398.195 ;
        END
    END p615
    PIN p616
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 398.405 208.355 398.475 ;
        END
    END p616
    PIN p617
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 402.045 208.355 402.115 ;
        END
    END p617
    PIN p618
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 402.325 208.355 402.395 ;
        END
    END p618
    PIN p619
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 405.965 208.355 406.035 ;
        END
    END p619
    PIN p620
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 406.245 208.355 406.315 ;
        END
    END p620
    PIN p621
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 409.885 208.355 409.955 ;
        END
    END p621
    PIN p622
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 410.165 208.355 410.235 ;
        END
    END p622
    PIN p623
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 413.805 208.355 413.875 ;
        END
    END p623
    PIN p624
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 414.085 208.355 414.155 ;
        END
    END p624
    PIN p625
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 417.725 208.355 417.795 ;
        END
    END p625
    PIN p626
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 418.005 208.355 418.075 ;
        END
    END p626
    PIN p627
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 421.645 208.355 421.715 ;
        END
    END p627
    PIN p628
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 421.925 208.355 421.995 ;
        END
    END p628
    PIN p629
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 425.565 208.355 425.635 ;
        END
    END p629
    PIN p630
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 425.845 208.355 425.915 ;
        END
    END p630
    PIN p631
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 429.485 208.355 429.555 ;
        END
    END p631
    PIN p632
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 429.765 208.355 429.835 ;
        END
    END p632
    PIN p633
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 433.405 208.355 433.475 ;
        END
    END p633
    PIN p634
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 433.685 208.355 433.755 ;
        END
    END p634
    PIN p635
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 437.325 208.355 437.395 ;
        END
    END p635
    PIN p636
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 437.605 208.355 437.675 ;
        END
    END p636
    PIN p637
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 441.245 208.355 441.315 ;
        END
    END p637
    PIN p638
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 441.525 208.355 441.595 ;
        END
    END p638
    PIN p639
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 445.165 208.355 445.235 ;
        END
    END p639
    PIN p640
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 445.445 208.355 445.515 ;
        END
    END p640
    PIN p641
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 449.085 208.355 449.155 ;
        END
    END p641
    PIN p642
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 449.365 208.355 449.435 ;
        END
    END p642
    PIN p643
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  208.285 453.005 208.355 453.075 ;
        END
    END p643
    PIN p644
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 425.845 162.995 425.915 ;
        END
    END p644
    PIN p645
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  162.925 429.485 162.995 429.555 ;
        END
    END p645
    PIN p646
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 343.245 717.395 343.315 ;
        END
    END p646
    PIN p647
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 343.525 717.395 343.595 ;
        END
    END p647
    PIN p648
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.885 347.445 717.955 347.515 ;
        END
    END p648
    PIN p649
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  703.885 374.605 703.955 374.675 ;
        END
    END p649
    PIN p650
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 374.885 717.395 374.955 ;
        END
    END p650
    PIN p651
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.885 375.165 717.955 375.235 ;
        END
    END p651
    PIN p652
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 378.525 717.395 378.595 ;
        END
    END p652
    PIN p653
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.885 378.805 717.955 378.875 ;
        END
    END p653
    PIN p654
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 355.285 717.395 355.355 ;
        END
    END p654
    PIN p655
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 358.925 717.395 358.995 ;
        END
    END p655
    PIN p656
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.325 359.205 717.395 359.275 ;
        END
    END p656
    PIN p657
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  717.885 363.125 717.955 363.195 ;
        END
    END p657
    PIN p658
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  708.365 327.565 708.435 327.635 ;
        END
    END p658
    OBS
      LAYER via2 ;
        RECT  0 0 838.04 661.92 ;
      LAYER metal2 ;
        RECT  0 0 838.04 661.92 ;
      LAYER via1 ;
        RECT  0 0 838.04 661.92 ;
      LAYER metal1 ;
        RECT  0 0 838.04 661.92 ;
    END
END fake_macro_newblue1_o330083

MACRO fake_macro_newblue1_o330084
    CLASS BLOCK ;
    SIZE 37.24 BY 99.12 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 10.325 1.715 10.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 8.925 33.075 8.995 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  19.565 8.085 19.635 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 10.045 1.715 10.115 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 38.045 1.715 38.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 16.485 1.715 16.555 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 18.165 1.715 18.235 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 19.845 1.715 19.915 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 21.525 1.715 21.595 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 23.205 1.715 23.275 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 24.885 1.715 24.955 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 26.565 1.715 26.635 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 28.245 1.715 28.315 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 29.925 1.715 29.995 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 31.605 1.715 31.675 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 33.285 1.715 33.355 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 34.965 1.715 35.035 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 36.645 1.715 36.715 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 38.325 1.715 38.395 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 40.005 1.715 40.075 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 41.685 1.715 41.755 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 43.365 1.715 43.435 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 45.045 1.715 45.115 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 46.725 1.715 46.795 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 48.405 1.715 48.475 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 50.085 1.715 50.155 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 51.765 1.715 51.835 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 53.445 1.715 53.515 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 55.125 1.715 55.195 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 56.805 1.715 56.875 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.485 1.715 58.555 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 61.845 1.715 61.915 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 63.525 1.715 63.595 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 65.205 1.715 65.275 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 66.885 1.715 66.955 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 68.565 1.715 68.635 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 70.245 1.715 70.315 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 71.925 1.715 71.995 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 73.605 1.715 73.675 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 75.285 1.715 75.355 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 76.965 1.715 77.035 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 78.645 1.715 78.715 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 80.325 1.715 80.395 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 82.005 1.715 82.075 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 82.005 35.315 82.075 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 80.325 35.315 80.395 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 78.645 35.315 78.715 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 76.965 35.315 77.035 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 75.285 35.315 75.355 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 73.605 35.315 73.675 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 71.925 35.315 71.995 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 70.245 35.315 70.315 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 68.565 35.315 68.635 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 66.885 35.315 66.955 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 65.205 35.315 65.275 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 63.525 35.315 63.595 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 61.845 35.315 61.915 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 60.165 35.315 60.235 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 58.485 35.315 58.555 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 56.805 35.315 56.875 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 55.125 35.315 55.195 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 53.445 35.315 53.515 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 51.765 35.315 51.835 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 50.085 35.315 50.155 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 48.405 35.315 48.475 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 46.725 35.315 46.795 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 45.045 35.315 45.115 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 43.365 35.315 43.435 ;
        END
    END p68
    PIN p69
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 41.685 35.315 41.755 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 40.005 35.315 40.075 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 38.325 35.315 38.395 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 36.645 35.315 36.715 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 34.965 35.315 35.035 ;
        END
    END p73
    PIN p74
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 33.285 35.315 33.355 ;
        END
    END p74
    PIN p75
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 31.605 35.315 31.675 ;
        END
    END p75
    PIN p76
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 29.925 35.315 29.995 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 28.245 35.315 28.315 ;
        END
    END p77
    PIN p78
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 26.565 35.315 26.635 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 24.885 35.315 24.955 ;
        END
    END p79
    PIN p80
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 23.205 35.315 23.275 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 21.525 35.315 21.595 ;
        END
    END p81
    PIN p82
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 19.845 35.315 19.915 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 18.165 35.315 18.235 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 16.485 35.315 16.555 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 9.485 34.755 9.555 ;
        END
    END p85
    OBS
      LAYER via2 ;
        RECT  0 0 37.24 99.12 ;
      LAYER metal2 ;
        RECT  0 0 37.24 99.12 ;
      LAYER via1 ;
        RECT  0 0 37.24 99.12 ;
      LAYER metal1 ;
        RECT  0 0 37.24 99.12 ;
    END
END fake_macro_newblue1_o330084

MACRO fake_macro_newblue1_o330180
    CLASS BLOCK ;
    SIZE 47.04 BY 38.64 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 12.845 27.475 12.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 15.925 10.115 15.995 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.765 15.925 16.835 15.995 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 15.925 10.675 15.995 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 29.925 11.235 29.995 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 29.925 11.795 29.995 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 29.925 10.115 29.995 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 29.925 25.795 29.995 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 29.925 9.555 29.995 ;
        END
    END p8
    OBS
      LAYER via2 ;
        RECT  0 0 47.04 38.64 ;
      LAYER metal2 ;
        RECT  0 0 47.04 38.64 ;
      LAYER via1 ;
        RECT  0 0 47.04 38.64 ;
      LAYER metal1 ;
        RECT  0 0 47.04 38.64 ;
    END
END fake_macro_newblue1_o330180

MACRO fake_macro_newblue1_o330181
    CLASS BLOCK ;
    SIZE 70 BY 82.32 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 66.325 22.435 66.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 66.325 29.155 66.395 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 66.325 58.275 66.395 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 60.725 61.635 60.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 59.325 61.635 59.395 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 61.005 61.635 61.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 82.005 61.635 82.075 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 61.285 61.635 61.355 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 60.445 61.635 60.515 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 55.685 61.635 55.755 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 52.045 61.635 52.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 55.965 61.635 56.035 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 52.325 61.635 52.395 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 20.405 61.635 20.475 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 15.645 61.635 15.715 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 15.365 61.635 15.435 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 25.725 61.635 25.795 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 32.725 61.635 32.795 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 26.845 61.635 26.915 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 17.045 61.635 17.115 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.125 15.645 62.195 15.715 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 20.685 61.635 20.755 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 57.365 61.635 57.435 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 20.965 61.635 21.035 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 46.165 61.635 46.235 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 50.925 61.635 50.995 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 45.885 61.635 45.955 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 32.165 61.635 32.235 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 51.205 61.635 51.275 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 47.285 61.635 47.355 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 30.485 61.635 30.555 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 27.125 61.635 27.195 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 22.085 61.635 22.155 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 34.405 61.635 34.475 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 30.765 61.635 30.835 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 32.445 61.635 32.515 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 35.245 61.635 35.315 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.125 30.765 62.195 30.835 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 23.765 61.635 23.835 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 59.045 61.635 59.115 ;
        END
    END p39
    OBS
      LAYER via2 ;
        RECT  0 0 70 82.32 ;
      LAYER metal2 ;
        RECT  0 0 70 82.32 ;
      LAYER via1 ;
        RECT  0 0 70 82.32 ;
      LAYER metal1 ;
        RECT  0 0 70 82.32 ;
    END
END fake_macro_newblue1_o330181

MACRO fake_macro_newblue1_o330182
    CLASS BLOCK ;
    SIZE 15.68 BY 157.92 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 78.085 14.035 78.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 80.885 14.035 80.955 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 83.685 1.715 83.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 81.725 1.715 81.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 73.045 14.035 73.115 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 81.445 14.035 81.515 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.125 1.155 76.195 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 71.925 1.155 71.995 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 79.205 14.035 79.275 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 83.405 1.715 83.475 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 33.565 14.035 33.635 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 27.685 14.035 27.755 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 23.765 14.035 23.835 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.045 14.035 10.115 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 8.085 14.035 8.155 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 4.165 14.035 4.235 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 29.645 14.035 29.715 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 13.965 14.035 14.035 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 19.845 14.035 19.915 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 62.965 14.035 63.035 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 49.245 14.035 49.315 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 39.445 14.035 39.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 66.885 14.035 66.955 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 53.165 14.035 53.235 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 43.365 14.035 43.435 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 70.805 14.035 70.875 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.085 14.035 57.155 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 47.285 14.035 47.355 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.885 14.035 115.955 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.965 14.035 112.035 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 100.205 14.035 100.275 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 86.765 14.035 86.835 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 92.365 14.035 92.435 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 119.805 14.035 119.875 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 106.365 14.035 106.435 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 102.445 14.035 102.515 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 96.285 14.035 96.355 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 145.565 14.035 145.635 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 133.805 14.035 133.875 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.045 14.035 122.115 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 151.165 14.035 151.235 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 139.405 14.035 139.475 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 125.965 14.035 126.035 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 153.405 14.035 153.475 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 141.645 14.035 141.715 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 131.565 14.035 131.635 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 65.765 14.035 65.835 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 69.685 14.035 69.755 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 142.485 14.035 142.555 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 146.405 14.035 146.475 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 150.325 14.035 150.395 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 154.245 14.035 154.315 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 111.405 1.715 111.475 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.885 14.035 3.955 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 84.525 14.035 84.595 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 2.485 14.035 2.555 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.405 14.035 6.475 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.325 14.035 10.395 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.245 14.035 14.315 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.165 14.035 18.235 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.085 14.035 22.155 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.005 14.035 26.075 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 29.925 14.035 29.995 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 33.845 14.035 33.915 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 37.765 14.035 37.835 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 41.685 14.035 41.755 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 45.605 14.035 45.675 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 49.525 14.035 49.595 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 53.445 14.035 53.515 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.365 14.035 57.435 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.285 14.035 61.355 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 65.205 14.035 65.275 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 69.125 14.035 69.195 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 88.165 14.035 88.235 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 92.085 14.035 92.155 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 96.005 14.035 96.075 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.925 14.035 99.995 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.845 14.035 103.915 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.765 14.035 107.835 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.685 14.035 111.755 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.605 14.035 115.675 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 119.525 14.035 119.595 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 123.445 14.035 123.515 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 127.365 14.035 127.435 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 131.285 14.035 131.355 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 135.205 14.035 135.275 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 139.125 14.035 139.195 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 143.045 14.035 143.115 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 146.965 14.035 147.035 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 150.885 14.035 150.955 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 154.805 14.035 154.875 ;
        END
    END p156
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 157.92 ;
      LAYER metal2 ;
        RECT  0 0 15.68 157.92 ;
      LAYER via1 ;
        RECT  0 0 15.68 157.92 ;
      LAYER metal1 ;
        RECT  0 0 15.68 157.92 ;
    END
END fake_macro_newblue1_o330182

MACRO fake_macro_newblue1_o330183
    CLASS BLOCK ;
    SIZE 15.68 BY 157.92 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.085 1.155 78.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 83.685 13.475 83.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.725 13.475 81.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 76.125 14.035 76.195 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 71.925 14.035 71.995 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.205 1.155 79.275 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 83.405 13.475 83.475 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 13.965 1.155 14.035 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.965 1.155 112.035 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.765 1.155 86.835 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.045 1.155 122.115 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.965 1.155 126.035 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 141.645 1.155 141.715 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 111.405 13.475 111.475 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.365 1.155 106.435 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 65.765 14.035 65.835 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 69.685 14.035 69.755 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 142.485 14.035 142.555 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 146.405 14.035 146.475 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 150.325 14.035 150.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 154.245 14.035 154.315 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p155
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 157.92 ;
      LAYER metal2 ;
        RECT  0 0 15.68 157.92 ;
      LAYER via1 ;
        RECT  0 0 15.68 157.92 ;
      LAYER metal1 ;
        RECT  0 0 15.68 157.92 ;
    END
END fake_macro_newblue1_o330183

MACRO fake_macro_newblue1_o330184
    CLASS BLOCK ;
    SIZE 15.68 BY 157.92 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.085 1.155 78.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 83.685 13.475 83.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.725 13.475 81.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 76.125 14.035 76.195 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 71.925 14.035 71.995 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.205 1.155 79.275 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 83.405 13.475 83.475 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.965 1.155 112.035 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.765 1.155 86.835 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.045 1.155 122.115 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.965 1.155 126.035 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 141.645 1.155 141.715 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 111.405 13.475 111.475 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.365 1.155 106.435 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 13.965 1.155 14.035 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 65.765 14.035 65.835 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 69.685 14.035 69.755 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 142.485 14.035 142.555 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 146.405 14.035 146.475 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 150.325 14.035 150.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 154.245 14.035 154.315 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p155
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 157.92 ;
      LAYER metal2 ;
        RECT  0 0 15.68 157.92 ;
      LAYER via1 ;
        RECT  0 0 15.68 157.92 ;
      LAYER metal1 ;
        RECT  0 0 15.68 157.92 ;
    END
END fake_macro_newblue1_o330184

MACRO fake_macro_newblue1_o330185
    CLASS BLOCK ;
    SIZE 15.68 BY 157.92 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 83.685 13.475 83.755 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.085 1.155 78.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.725 13.475 81.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 76.125 14.035 76.195 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 71.925 14.035 71.995 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.205 1.155 79.275 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 83.405 13.475 83.475 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.965 1.155 112.035 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.765 1.155 86.835 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.045 1.155 122.115 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 141.645 1.155 141.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.965 1.155 126.035 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 111.405 13.475 111.475 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.365 1.155 106.435 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 13.965 1.155 14.035 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 65.765 14.035 65.835 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 69.685 14.035 69.755 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 142.485 14.035 142.555 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 146.405 14.035 146.475 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 150.325 14.035 150.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 154.245 14.035 154.315 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p155
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 157.92 ;
      LAYER metal2 ;
        RECT  0 0 15.68 157.92 ;
      LAYER via1 ;
        RECT  0 0 15.68 157.92 ;
      LAYER metal1 ;
        RECT  0 0 15.68 157.92 ;
    END
END fake_macro_newblue1_o330185

MACRO fake_macro_newblue1_o330186
    CLASS BLOCK ;
    SIZE 39.2 BY 157.92 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 81.725 36.995 81.795 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 76.125 37.555 76.195 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 71.925 37.555 71.995 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.085 1.155 78.155 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.205 1.155 79.275 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 78.085 1.715 78.155 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 79.205 1.715 79.275 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 78.085 3.395 78.155 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 79.205 3.395 79.275 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 83.685 36.995 83.755 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 83.405 36.995 83.475 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 13.965 1.155 14.035 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.125 1.155 6.195 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.805 1.155 21.875 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 68.845 1.155 68.915 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.005 1.155 61.075 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 114.205 1.155 114.275 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.285 1.155 110.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 94.605 1.155 94.675 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.685 1.155 90.755 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.485 1.155 135.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.885 1.155 129.955 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.645 1.155 127.715 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.045 1.155 122.115 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.085 1.155 155.155 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 149.485 1.155 149.555 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.245 1.155 147.315 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 141.645 1.155 141.715 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 111.405 36.995 111.475 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 3.045 37.555 3.115 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 6.965 37.555 7.035 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 10.885 37.555 10.955 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 14.805 37.555 14.875 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 18.725 37.555 18.795 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 22.645 37.555 22.715 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 26.565 37.555 26.635 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 30.485 37.555 30.555 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 34.405 37.555 34.475 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 38.325 37.555 38.395 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 42.245 37.555 42.315 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 46.165 37.555 46.235 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 50.085 37.555 50.155 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 54.005 37.555 54.075 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 57.925 37.555 57.995 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 61.845 37.555 61.915 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 65.765 37.555 65.835 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 69.685 37.555 69.755 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 87.605 37.555 87.675 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 91.525 37.555 91.595 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 95.445 37.555 95.515 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 99.365 37.555 99.435 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 103.285 37.555 103.355 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 107.205 37.555 107.275 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 111.125 37.555 111.195 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 115.045 37.555 115.115 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 118.965 37.555 119.035 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 122.885 37.555 122.955 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 126.805 37.555 126.875 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 130.725 37.555 130.795 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 134.645 37.555 134.715 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 138.565 37.555 138.635 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 142.485 37.555 142.555 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 146.405 37.555 146.475 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 150.325 37.555 150.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 154.245 37.555 154.315 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p159
    OBS
      LAYER via2 ;
        RECT  0 0 39.2 157.92 ;
      LAYER metal2 ;
        RECT  0 0 39.2 157.92 ;
      LAYER via1 ;
        RECT  0 0 39.2 157.92 ;
      LAYER metal1 ;
        RECT  0 0 39.2 157.92 ;
    END
END fake_macro_newblue1_o330186

MACRO fake_macro_newblue1_o330227
    CLASS BLOCK ;
    SIZE 39.2 BY 268.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 138.565 36.995 138.635 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.245 1.155 252.315 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.165 1.155 256.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.085 1.155 260.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.005 1.155 264.075 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.125 1.155 6.195 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.645 1.155 78.715 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 98.245 1.155 98.315 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.765 1.155 121.835 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.245 1.155 147.315 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 149.485 1.155 149.555 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.925 1.155 162.995 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.765 1.155 170.835 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.605 1.155 178.675 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.285 1.155 194.355 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.125 1.155 202.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.965 1.155 210.035 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 212.205 1.155 212.275 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.805 1.155 217.875 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.645 1.155 225.715 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.485 1.155 233.555 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.325 1.155 241.395 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 243.565 1.155 243.635 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 249.165 1.155 249.235 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 251.405 1.155 251.475 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.005 1.155 257.075 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.925 1.155 260.995 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.845 1.155 264.915 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 131.005 37.555 131.075 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 126.805 37.555 126.875 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.965 1.155 133.035 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 132.965 1.715 133.035 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 132.965 3.395 133.035 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 136.605 36.995 136.675 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.325 1.155 136.395 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.085 1.155 134.155 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 134.085 1.715 134.155 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 134.085 3.395 134.155 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 138.285 36.995 138.355 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 166.285 36.995 166.355 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 3.045 37.555 3.115 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 6.965 37.555 7.035 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 10.885 37.555 10.955 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 14.805 37.555 14.875 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 18.725 37.555 18.795 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 22.645 37.555 22.715 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 26.565 37.555 26.635 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 30.485 37.555 30.555 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 34.405 37.555 34.475 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 38.325 37.555 38.395 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 42.245 37.555 42.315 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 46.165 37.555 46.235 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 50.085 37.555 50.155 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 54.005 37.555 54.075 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 57.925 37.555 57.995 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 61.845 37.555 61.915 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 65.765 37.555 65.835 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 69.685 37.555 69.755 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 73.605 37.555 73.675 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 77.525 37.555 77.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 81.445 37.555 81.515 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 85.365 37.555 85.435 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 89.285 37.555 89.355 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 93.205 37.555 93.275 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 97.125 37.555 97.195 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 101.045 37.555 101.115 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 104.965 37.555 105.035 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 108.885 37.555 108.955 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 112.805 37.555 112.875 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 116.725 37.555 116.795 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 120.645 37.555 120.715 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 124.565 37.555 124.635 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 142.485 37.555 142.555 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 146.405 37.555 146.475 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 150.325 37.555 150.395 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 154.245 37.555 154.315 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 158.165 37.555 158.235 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 162.085 37.555 162.155 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 166.005 37.555 166.075 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 169.925 37.555 169.995 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 173.845 37.555 173.915 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 177.765 37.555 177.835 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 181.685 37.555 181.755 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 185.605 37.555 185.675 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 189.525 37.555 189.595 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 193.445 37.555 193.515 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 197.365 37.555 197.435 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 201.285 37.555 201.355 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 205.205 37.555 205.275 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 209.125 37.555 209.195 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 213.045 37.555 213.115 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 216.965 37.555 217.035 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 220.885 37.555 220.955 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 224.805 37.555 224.875 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 228.725 37.555 228.795 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 232.645 37.555 232.715 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 236.565 37.555 236.635 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 240.485 37.555 240.555 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 244.405 37.555 244.475 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 248.325 37.555 248.395 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 252.245 37.555 252.315 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 256.165 37.555 256.235 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 260.085 37.555 260.155 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 264.005 37.555 264.075 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.805 1.155 252.875 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.645 1.155 260.715 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p271
    OBS
      LAYER via2 ;
        RECT  0 0 39.2 268.8 ;
      LAYER metal2 ;
        RECT  0 0 39.2 268.8 ;
      LAYER via1 ;
        RECT  0 0 39.2 268.8 ;
      LAYER metal1 ;
        RECT  0 0 39.2 268.8 ;
    END
END fake_macro_newblue1_o330227

MACRO fake_macro_newblue1_o330228
    CLASS BLOCK ;
    SIZE 11.76 BY 268.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 264.565 10.115 264.635 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 138.565 1.715 138.635 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 120.645 10.115 120.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 124.565 10.115 124.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 252.245 10.115 252.315 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 256.165 10.115 256.235 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 260.085 10.115 260.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 264.005 10.115 264.075 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 2.205 10.115 2.275 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 8.085 10.115 8.155 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 12.005 10.115 12.075 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 15.925 10.115 15.995 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 19.845 10.115 19.915 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 23.765 10.115 23.835 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 27.685 10.115 27.755 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 31.605 10.115 31.675 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 35.525 10.115 35.595 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 37.485 10.115 37.555 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 43.365 10.115 43.435 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 45.325 10.115 45.395 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 51.205 10.115 51.275 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 53.165 10.115 53.235 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 59.045 10.115 59.115 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.005 10.115 61.075 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 66.885 10.115 66.955 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 70.805 10.115 70.875 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 74.725 10.115 74.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 78.645 10.115 78.715 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 82.565 10.115 82.635 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 86.485 10.115 86.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 90.405 10.115 90.475 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 94.325 10.115 94.395 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 96.285 10.115 96.355 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 102.165 10.115 102.235 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.125 10.115 104.195 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 110.005 10.115 110.075 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 111.965 10.115 112.035 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 117.845 10.115 117.915 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 119.805 10.115 119.875 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 125.685 10.115 125.755 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 143.325 10.115 143.395 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 145.565 10.115 145.635 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 151.165 10.115 151.235 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 155.085 10.115 155.155 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 159.005 10.115 159.075 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.925 10.115 162.995 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.845 10.115 166.915 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 170.765 10.115 170.835 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 174.685 10.115 174.755 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 178.605 10.115 178.675 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 182.525 10.115 182.595 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 186.445 10.115 186.515 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 188.685 10.115 188.755 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 194.285 10.115 194.355 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 196.525 10.115 196.595 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 202.125 10.115 202.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 204.365 10.115 204.435 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.965 10.115 210.035 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.885 10.115 213.955 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 217.805 10.115 217.875 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 221.725 10.115 221.795 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 225.645 10.115 225.715 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 229.565 10.115 229.635 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 233.485 10.115 233.555 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 237.405 10.115 237.475 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 241.325 10.115 241.395 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 245.245 10.115 245.315 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 247.485 10.115 247.555 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 253.085 10.115 253.155 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 255.325 10.115 255.395 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 260.925 10.115 260.995 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 263.165 10.115 263.235 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 127.925 10.115 127.995 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.005 1.155 131.075 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 139.405 10.115 139.475 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 136.605 1.715 136.675 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 136.325 10.115 136.395 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 135.765 10.115 135.835 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 138.285 1.715 138.355 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 166.285 1.715 166.355 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.245 1.155 252.315 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.165 1.155 256.235 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.085 1.155 260.155 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.005 1.155 264.075 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 2.485 10.115 2.555 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.405 10.115 6.475 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.325 10.115 10.395 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.245 10.115 14.315 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.165 10.115 18.235 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.085 10.115 22.155 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.005 10.115 26.075 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 29.925 10.115 29.995 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 33.845 10.115 33.915 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 37.765 10.115 37.835 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 41.685 10.115 41.755 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 45.605 10.115 45.675 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 49.525 10.115 49.595 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 53.445 10.115 53.515 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.365 10.115 57.435 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.285 10.115 61.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.205 10.115 65.275 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.125 10.115 69.195 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.045 10.115 73.115 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 76.965 10.115 77.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 80.885 10.115 80.955 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 84.805 10.115 84.875 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 88.725 10.115 88.795 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 92.645 10.115 92.715 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 96.565 10.115 96.635 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 100.485 10.115 100.555 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.405 10.115 104.475 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.325 10.115 108.395 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.245 10.115 112.315 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.165 10.115 116.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 120.085 10.115 120.155 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 124.005 10.115 124.075 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 143.045 10.115 143.115 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.965 10.115 147.035 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.885 10.115 150.955 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.805 10.115 154.875 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.725 10.115 158.795 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.645 10.115 162.715 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.565 10.115 166.635 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 170.485 10.115 170.555 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 174.405 10.115 174.475 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 178.325 10.115 178.395 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 182.245 10.115 182.315 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 186.165 10.115 186.235 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 190.085 10.115 190.155 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 194.005 10.115 194.075 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.925 10.115 197.995 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.845 10.115 201.915 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.765 10.115 205.835 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.685 10.115 209.755 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.605 10.115 213.675 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 217.525 10.115 217.595 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 221.445 10.115 221.515 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 225.365 10.115 225.435 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 229.285 10.115 229.355 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 233.205 10.115 233.275 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 237.125 10.115 237.195 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 241.045 10.115 241.115 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.965 10.115 245.035 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.885 10.115 248.955 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 252.805 10.115 252.875 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 256.725 10.115 256.795 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 260.645 10.115 260.715 ;
        END
    END p265
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER via1 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal1 ;
        RECT  0 0 11.76 268.8 ;
    END
END fake_macro_newblue1_o330228

MACRO fake_macro_newblue1_o330273
    CLASS BLOCK ;
    SIZE 103.88 BY 131.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 20.125 10.675 20.195 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.205 1.645 100.275 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 1.645 98.595 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  92.365 1.645 92.435 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 1.645 90.755 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.885 1.645 87.955 1.715 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 1.645 86.275 1.715 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  84.525 1.645 84.595 1.715 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 1.645 82.915 1.715 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 1.645 80.675 1.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 1.645 78.995 1.715 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.245 1.645 77.315 1.715 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 1.645 75.635 1.715 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 1.645 69.475 1.715 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 1.645 67.795 1.715 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 1.645 65.555 1.715 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 1.645 63.875 1.715 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.125 1.645 62.195 1.715 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 1.645 60.515 1.715 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 1.645 58.275 1.715 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 1.645 56.595 1.715 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.725 1.645 53.795 1.715 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 1.645 52.115 1.715 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 1.645 50.435 1.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 1.645 48.755 1.715 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  46.445 1.645 46.515 1.715 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 1.645 44.835 1.715 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 1.645 43.155 1.715 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 1.645 41.475 1.715 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 1.645 35.315 1.715 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 1.645 33.635 1.715 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.325 1.645 31.395 1.715 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 1.645 29.715 1.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 1.645 28.035 1.715 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 1.645 26.355 1.715 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.045 1.645 24.115 1.715 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 1.645 22.435 1.715 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 24.605 3.955 24.675 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 26.845 3.955 26.915 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 54.565 3.955 54.635 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 29.085 3.955 29.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 29.365 4.515 29.435 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 31.325 3.955 31.395 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 20.125 3.955 20.195 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 22.365 3.955 22.435 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.325 1.645 101.395 1.715 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 1.645 99.155 1.715 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 1.645 93.555 1.715 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 1.645 91.315 1.715 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 1.645 89.075 1.715 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 1.645 86.835 1.715 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 1.645 85.155 1.715 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 1.645 83.475 1.715 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 1.645 81.795 1.715 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 1.645 79.555 1.715 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.645 77.875 1.715 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 1.645 76.195 1.715 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 1.645 70.035 1.715 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 1.645 68.355 1.715 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 1.645 66.675 1.715 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 1.645 64.435 1.715 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 1.645 62.755 1.715 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 1.645 61.075 1.715 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 1.645 59.395 1.715 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.645 57.155 1.715 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 1.645 54.915 1.715 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 1.645 52.675 1.715 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 1.645 50.995 1.715 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 1.645 49.315 1.715 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 1.645 47.635 1.715 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 1.645 45.395 1.715 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 1.645 43.715 1.715 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 1.645 42.035 1.715 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 1.645 35.875 1.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 1.645 34.195 1.715 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 1.645 32.515 1.715 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 1.645 30.275 1.715 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 1.645 28.595 1.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 1.645 26.915 1.715 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 1.645 25.235 1.715 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 1.645 22.995 1.715 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 12.005 3.955 12.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 31.605 4.515 31.675 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 12.845 12.915 12.915 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 5.565 12.355 5.635 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 1.925 11.795 1.995 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.925 6.755 1.995 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 6.405 7.875 6.475 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 6.685 5.635 6.755 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 13.125 2.275 13.195 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 5.565 16.275 5.635 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 5.565 14.595 5.635 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.085 5.565 15.155 5.635 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 33.285 12.355 33.355 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 22.645 4.515 22.715 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 20.125 3.395 20.195 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 20.405 4.515 20.475 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 17.885 3.395 17.955 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 17.885 3.955 17.955 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 31.325 3.395 31.395 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 31.045 4.515 31.115 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 29.085 3.395 29.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 28.805 4.515 28.875 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 26.845 3.395 26.915 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 27.125 4.515 27.195 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 24.605 3.395 24.675 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 24.885 4.515 24.955 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 22.365 3.395 22.435 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 12.005 3.395 12.075 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 13.405 2.275 13.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 18.165 23.555 18.235 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 18.165 25.235 18.235 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 18.165 27.475 18.235 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 18.165 29.155 18.235 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 18.165 30.835 18.235 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 18.165 32.515 18.235 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 18.165 34.755 18.235 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 18.165 36.435 18.235 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 18.165 42.595 18.235 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 18.165 44.275 18.235 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 18.165 45.955 18.235 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 18.165 47.635 18.235 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 18.165 49.875 18.235 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 18.165 51.555 18.235 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 18.165 53.235 18.235 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 18.165 54.915 18.235 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 18.165 57.715 18.235 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 18.165 59.395 18.235 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 18.165 61.635 18.235 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.245 18.165 63.315 18.235 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 18.165 64.995 18.235 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 18.165 66.675 18.235 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 18.165 68.915 18.235 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 18.165 70.595 18.235 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 18.165 76.755 18.235 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.365 18.165 78.435 18.235 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 18.165 80.115 18.235 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 18.165 81.795 18.235 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 18.165 84.035 18.235 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.645 18.165 85.715 18.235 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 18.165 87.395 18.235 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 18.165 89.075 18.235 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 18.165 91.875 18.235 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 18.165 93.555 18.235 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.645 18.165 99.715 18.235 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.325 18.165 101.395 18.235 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 41.125 2.275 41.195 ;
        END
    END p146
    OBS
      LAYER via2 ;
        RECT  0 0 104.02 131.04 ;
      LAYER metal2 ;
        RECT  0 0 104.02 131.04 ;
      LAYER via1 ;
        RECT  0 0 104.02 131.04 ;
      LAYER metal1 ;
        RECT  0 0 104.02 131.04 ;
    END
END fake_macro_newblue1_o330273

MACRO fake_macro_newblue1_o330274
    CLASS BLOCK ;
    SIZE 168.56 BY 99.12 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  165.165 97.125 165.235 97.195 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.005 97.125 159.075 97.195 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  156.205 97.125 156.275 97.195 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  154.525 97.125 154.595 97.195 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.845 97.125 152.915 97.195 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.165 97.125 151.235 97.195 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.925 97.125 148.995 97.195 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.245 97.125 147.315 97.195 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.565 97.125 145.635 97.195 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  143.885 97.125 143.955 97.195 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.725 97.125 137.795 97.195 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 97.125 136.115 97.195 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.805 97.125 133.875 97.195 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.125 97.125 132.195 97.195 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  130.445 97.125 130.515 97.195 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  128.765 97.125 128.835 97.195 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  126.525 97.125 126.595 97.195 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  124.845 97.125 124.915 97.195 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 97.125 122.115 97.195 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 97.125 120.435 97.195 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.685 97.125 118.755 97.195 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 97.125 117.075 97.195 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.765 97.125 114.835 97.195 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.085 97.125 113.155 97.195 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  111.405 97.125 111.475 97.195 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  109.725 97.125 109.795 97.195 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.565 97.125 103.635 97.195 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.885 97.125 101.955 97.195 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.645 97.125 99.715 97.195 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.965 97.125 98.035 97.195 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 97.125 96.355 97.195 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 97.125 94.675 97.195 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  92.365 97.125 92.435 97.195 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 97.125 90.755 97.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.885 97.125 87.955 97.195 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 97.125 86.275 97.195 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  84.525 97.125 84.595 97.195 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 97.125 82.915 97.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 97.125 80.675 97.195 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 97.125 78.995 97.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.245 97.125 77.315 97.195 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 97.125 75.635 97.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 97.125 69.475 97.195 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 97.125 67.795 97.195 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 97.125 65.555 97.195 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 97.125 63.875 97.195 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.125 97.125 62.195 97.195 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 97.125 60.515 97.195 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 97.125 58.275 97.195 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 97.125 56.595 97.195 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.725 97.125 53.795 97.195 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 97.125 52.115 97.195 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 97.125 50.435 97.195 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 97.125 48.755 97.195 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  46.445 97.125 46.515 97.195 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 97.125 44.835 97.195 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 97.125 43.155 97.195 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 97.125 41.475 97.195 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 97.125 35.315 97.195 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 97.125 33.635 97.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.325 97.125 31.395 97.195 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 97.125 29.715 97.195 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 97.125 28.035 97.195 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 97.125 26.355 97.195 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.045 97.125 24.115 97.195 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 97.125 22.435 97.195 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 93.205 12.355 93.275 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 96.845 6.755 96.915 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 93.205 16.275 93.275 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.085 93.205 15.155 93.275 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 98.805 12.355 98.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 86.765 3.395 86.835 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 76.405 3.955 76.475 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 78.645 3.955 78.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 67.445 3.955 67.515 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 95.165 3.955 95.235 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 69.685 3.955 69.755 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 69.965 4.515 70.035 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 71.925 3.955 71.995 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 72.205 4.515 72.275 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 85.925 12.915 85.995 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 97.125 22.995 97.195 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 97.125 25.235 97.195 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 97.125 26.915 97.195 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 97.125 28.595 97.195 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 97.125 30.275 97.195 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 97.125 32.515 97.195 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 97.125 34.195 97.195 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 97.125 35.875 97.195 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 97.125 42.035 97.195 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 97.125 43.715 97.195 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 97.125 45.395 97.195 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 97.125 47.635 97.195 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 97.125 49.315 97.195 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 97.125 50.995 97.195 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 97.125 52.675 97.195 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 97.125 54.915 97.195 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 97.125 57.155 97.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 97.125 59.395 97.195 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 97.125 61.075 97.195 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 97.125 62.755 97.195 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 97.125 64.435 97.195 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 97.125 66.675 97.195 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 97.125 68.355 97.195 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 97.125 70.035 97.195 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 97.125 76.195 97.195 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 97.125 77.875 97.195 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 97.125 79.555 97.195 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 97.125 81.795 97.195 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 97.125 83.475 97.195 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 97.125 85.155 97.195 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 97.125 86.835 97.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 97.125 89.075 97.195 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 97.125 91.315 97.195 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 97.125 93.555 97.195 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 97.125 95.235 97.195 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 97.125 96.915 97.195 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 97.125 98.595 97.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 97.125 100.835 97.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 97.125 102.515 97.195 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.125 97.125 104.195 97.195 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.285 97.125 110.355 97.195 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  111.965 97.125 112.035 97.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.645 97.125 113.715 97.195 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  115.885 97.125 115.955 97.195 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.565 97.125 117.635 97.195 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.245 97.125 119.315 97.195 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 97.125 120.995 97.195 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  123.165 97.125 123.235 97.195 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.405 97.125 125.475 97.195 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  127.645 97.125 127.715 97.195 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.325 97.125 129.395 97.195 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  131.005 97.125 131.075 97.195 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.685 97.125 132.755 97.195 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.925 97.125 134.995 97.195 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.605 97.125 136.675 97.195 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  138.285 97.125 138.355 97.195 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  144.445 97.125 144.515 97.195 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  146.125 97.125 146.195 97.195 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.805 97.125 147.875 97.195 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  150.045 97.125 150.115 97.195 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.725 97.125 151.795 97.195 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  153.405 97.125 153.475 97.195 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.085 97.125 155.155 97.195 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  157.325 97.125 157.395 97.195 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 97.125 159.635 97.195 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  165.725 97.125 165.795 97.195 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 96.845 11.795 96.915 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 92.365 7.875 92.435 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 92.085 5.635 92.155 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 85.645 2.275 85.715 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 93.205 14.595 93.275 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 76.685 4.515 76.755 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 78.645 3.395 78.715 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 78.925 4.515 78.995 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 80.885 3.395 80.955 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 80.885 3.955 80.955 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 67.445 3.395 67.515 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 67.725 4.515 67.795 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 69.685 3.395 69.755 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 69.405 4.515 69.475 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 71.925 3.395 71.995 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 71.645 4.515 71.715 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 74.165 3.395 74.235 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 74.165 3.955 74.235 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 76.405 3.395 76.475 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 86.765 3.955 86.835 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 85.365 2.275 85.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 80.605 23.555 80.675 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 80.605 25.235 80.675 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 80.605 27.475 80.675 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 80.605 29.155 80.675 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 80.605 30.835 80.675 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 80.605 32.515 80.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 80.605 34.755 80.675 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 80.605 36.435 80.675 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 80.605 42.595 80.675 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 80.605 44.275 80.675 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 80.605 45.955 80.675 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 80.605 47.635 80.675 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 80.605 49.875 80.675 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 80.605 51.555 80.675 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 80.605 53.235 80.675 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 80.605 54.915 80.675 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 80.605 57.715 80.675 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 80.605 59.395 80.675 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 80.605 61.635 80.675 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.245 80.605 63.315 80.675 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 80.605 64.995 80.675 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 80.605 66.675 80.675 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 80.605 68.915 80.675 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 80.605 70.595 80.675 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 80.605 76.755 80.675 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.365 80.605 78.435 80.675 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 80.605 80.115 80.675 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 80.605 81.795 80.675 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 80.605 84.035 80.675 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.645 80.605 85.715 80.675 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 80.605 87.395 80.675 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 80.605 89.075 80.675 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 80.605 91.875 80.675 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 80.605 93.555 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 80.605 95.795 80.675 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 80.605 97.475 80.675 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 80.605 99.155 80.675 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 80.605 100.835 80.675 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 80.605 103.075 80.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.685 80.605 104.755 80.675 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.845 80.605 110.915 80.675 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  112.525 80.605 112.595 80.675 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.205 80.605 114.275 80.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  115.885 80.605 115.955 80.675 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.125 80.605 118.195 80.675 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 80.605 119.875 80.675 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 80.605 121.555 80.675 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  123.165 80.605 123.235 80.675 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 80.605 126.035 80.675 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  127.645 80.605 127.715 80.675 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.885 80.605 129.955 80.675 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  131.565 80.605 131.635 80.675 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 80.605 133.315 80.675 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.925 80.605 134.995 80.675 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.165 80.605 137.235 80.675 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  138.845 80.605 138.915 80.675 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.005 80.605 145.075 80.675 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  146.685 80.605 146.755 80.675 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.365 80.605 148.435 80.675 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  150.045 80.605 150.115 80.675 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.285 80.605 152.355 80.675 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  153.965 80.605 154.035 80.675 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.645 80.605 155.715 80.675 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  157.325 80.605 157.395 80.675 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.125 80.605 160.195 80.675 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  166.285 80.605 166.355 80.675 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 98.805 2.275 98.875 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 78.645 10.675 78.715 ;
        END
    END p235
    OBS
      LAYER via2 ;
        RECT  0 0 168.7 99.12 ;
      LAYER metal2 ;
        RECT  0 0 168.7 99.12 ;
      LAYER via1 ;
        RECT  0 0 168.7 99.12 ;
      LAYER metal1 ;
        RECT  0 0 168.7 99.12 ;
    END
END fake_macro_newblue1_o330274

MACRO fake_macro_newblue1_o330275
    CLASS BLOCK ;
    SIZE 168.56 BY 99.12 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 78.645 10.675 78.715 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 93.205 12.355 93.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 96.845 6.755 96.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 93.205 16.275 93.275 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.085 93.205 15.155 93.275 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 98.805 12.355 98.875 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 86.765 3.395 86.835 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 96.845 11.795 96.915 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 92.365 7.875 92.435 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 85.645 2.275 85.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 93.205 14.595 93.275 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 76.405 3.955 76.475 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 78.645 3.395 78.715 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 78.645 3.955 78.715 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 80.885 3.395 80.955 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 80.885 3.955 80.955 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 67.445 3.395 67.515 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 67.445 3.955 67.515 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 69.685 3.395 69.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 69.685 3.955 69.755 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 71.925 3.395 71.995 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 71.925 3.955 71.995 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 74.165 3.395 74.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 74.165 3.955 74.235 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 76.405 3.395 76.475 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 98.805 3.955 98.875 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 78.925 4.515 78.995 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 67.725 4.515 67.795 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 67.165 4.515 67.235 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 69.965 4.515 70.035 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 69.405 4.515 69.475 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 72.205 4.515 72.275 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 71.645 4.515 71.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  109.725 97.125 109.795 97.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 97.125 96.355 97.195 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 97.125 86.275 97.195 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.245 97.125 77.315 97.195 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 97.125 63.875 97.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.725 97.125 53.795 97.195 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 97.125 44.835 97.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.325 97.125 31.395 97.195 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 97.125 22.435 97.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.845 97.125 152.915 97.195 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  143.885 97.125 143.955 97.195 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  130.445 97.125 130.515 97.195 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 97.125 120.435 97.195 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  111.405 97.125 111.475 97.195 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.965 97.125 98.035 97.195 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.885 97.125 87.955 97.195 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 97.125 78.995 97.195 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 97.125 65.555 97.195 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 97.125 56.595 97.195 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  46.445 97.125 46.515 97.195 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 97.125 33.635 97.195 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.045 97.125 24.115 97.195 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.005 97.125 159.075 97.195 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  156.205 97.125 156.275 97.195 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  154.525 97.125 154.595 97.195 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.925 97.125 148.995 97.195 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.565 97.125 145.635 97.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.725 97.125 137.795 97.195 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 97.125 136.115 97.195 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.125 97.125 132.195 97.195 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 97.125 122.115 97.195 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 97.125 117.075 97.195 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.765 97.125 114.835 97.195 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.885 97.125 101.955 97.195 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  92.365 97.125 92.435 97.195 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 97.125 69.475 97.195 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 97.125 60.515 97.195 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 97.125 52.115 97.195 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 97.125 26.355 97.195 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.245 97.125 147.315 97.195 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.805 97.125 133.875 97.195 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.565 97.125 103.635 97.195 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  84.525 97.125 84.595 97.195 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 97.125 67.795 97.195 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 97.125 48.755 97.195 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 97.125 41.475 97.195 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 97.125 29.715 97.195 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 97.125 28.035 97.195 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.165 97.125 151.235 97.195 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  128.765 97.125 128.835 97.195 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  126.525 97.125 126.595 97.195 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  124.845 97.125 124.915 97.195 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.685 97.125 118.755 97.195 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.645 97.125 99.715 97.195 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 97.125 94.675 97.195 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 97.125 90.755 97.195 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 97.125 82.915 97.195 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 97.125 80.675 97.195 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 97.125 75.635 97.195 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.125 97.125 62.195 97.195 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 97.125 58.275 97.195 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 97.125 50.435 97.195 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 97.125 43.155 97.195 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 97.125 35.315 97.195 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  165.165 97.125 165.235 97.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.085 97.125 113.155 97.195 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 85.925 12.915 85.995 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 97.125 22.995 97.195 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 97.125 25.235 97.195 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 97.125 26.915 97.195 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 97.125 28.595 97.195 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 97.125 30.275 97.195 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 97.125 32.515 97.195 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 97.125 34.195 97.195 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 97.125 35.875 97.195 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 97.125 42.035 97.195 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 97.125 43.715 97.195 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 97.125 45.395 97.195 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 97.125 47.635 97.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 97.125 49.315 97.195 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 97.125 50.995 97.195 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 97.125 52.675 97.195 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 97.125 54.915 97.195 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 97.125 57.155 97.195 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 97.125 59.395 97.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 97.125 61.075 97.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 97.125 62.755 97.195 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 97.125 64.435 97.195 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 97.125 66.675 97.195 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 97.125 68.355 97.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 97.125 70.035 97.195 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 97.125 76.195 97.195 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 97.125 77.875 97.195 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 97.125 79.555 97.195 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 97.125 81.795 97.195 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 97.125 83.475 97.195 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 97.125 85.155 97.195 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 97.125 86.835 97.195 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 97.125 89.075 97.195 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 97.125 91.315 97.195 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 97.125 93.555 97.195 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 97.125 95.235 97.195 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 97.125 96.915 97.195 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 97.125 98.595 97.195 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 97.125 100.835 97.195 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 97.125 102.515 97.195 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.125 97.125 104.195 97.195 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.285 97.125 110.355 97.195 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  111.965 97.125 112.035 97.195 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.645 97.125 113.715 97.195 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  115.885 97.125 115.955 97.195 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.565 97.125 117.635 97.195 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.245 97.125 119.315 97.195 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 97.125 120.995 97.195 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  123.165 97.125 123.235 97.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.405 97.125 125.475 97.195 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  127.645 97.125 127.715 97.195 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.325 97.125 129.395 97.195 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  131.005 97.125 131.075 97.195 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.685 97.125 132.755 97.195 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.925 97.125 134.995 97.195 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.605 97.125 136.675 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  138.285 97.125 138.355 97.195 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  144.445 97.125 144.515 97.195 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  146.125 97.125 146.195 97.195 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.805 97.125 147.875 97.195 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  150.045 97.125 150.115 97.195 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.725 97.125 151.795 97.195 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  153.405 97.125 153.475 97.195 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.085 97.125 155.155 97.195 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  157.325 97.125 157.395 97.195 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 97.125 159.635 97.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  165.725 97.125 165.795 97.195 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 92.085 5.635 92.155 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 86.765 3.955 86.835 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 85.365 2.275 85.435 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 80.605 23.555 80.675 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 80.605 25.235 80.675 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 80.605 27.475 80.675 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 80.605 29.155 80.675 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 80.605 30.835 80.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 80.605 32.515 80.675 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 80.605 34.755 80.675 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 80.605 36.435 80.675 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 80.605 42.595 80.675 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 80.605 44.275 80.675 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 80.605 45.955 80.675 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 80.605 47.635 80.675 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 80.605 49.875 80.675 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 80.605 51.555 80.675 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 80.605 53.235 80.675 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 80.605 54.915 80.675 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 80.605 57.715 80.675 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 80.605 59.395 80.675 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 80.605 61.635 80.675 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.245 80.605 63.315 80.675 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 80.605 64.995 80.675 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 80.605 66.675 80.675 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 80.605 68.915 80.675 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 80.605 70.595 80.675 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 80.605 76.755 80.675 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.365 80.605 78.435 80.675 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 80.605 80.115 80.675 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 80.605 81.795 80.675 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 80.605 84.035 80.675 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.645 80.605 85.715 80.675 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 80.605 87.395 80.675 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 80.605 89.075 80.675 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 80.605 91.875 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 80.605 93.555 80.675 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 80.605 95.795 80.675 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 80.605 97.475 80.675 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 80.605 99.155 80.675 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 80.605 100.835 80.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 80.605 103.075 80.675 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.685 80.605 104.755 80.675 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.845 80.605 110.915 80.675 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  112.525 80.605 112.595 80.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.205 80.605 114.275 80.675 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  115.885 80.605 115.955 80.675 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.125 80.605 118.195 80.675 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 80.605 119.875 80.675 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 80.605 121.555 80.675 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  123.165 80.605 123.235 80.675 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 80.605 126.035 80.675 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  127.645 80.605 127.715 80.675 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.885 80.605 129.955 80.675 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  131.565 80.605 131.635 80.675 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 80.605 133.315 80.675 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.925 80.605 134.995 80.675 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.165 80.605 137.235 80.675 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  138.845 80.605 138.915 80.675 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.005 80.605 145.075 80.675 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  146.685 80.605 146.755 80.675 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.365 80.605 148.435 80.675 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  150.045 80.605 150.115 80.675 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.285 80.605 152.355 80.675 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  153.965 80.605 154.035 80.675 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.645 80.605 155.715 80.675 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  157.325 80.605 157.395 80.675 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.125 80.605 160.195 80.675 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  166.285 80.605 166.355 80.675 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 98.805 2.275 98.875 ;
        END
    END p235
    OBS
      LAYER via2 ;
        RECT  0 0 168.7 99.12 ;
      LAYER metal2 ;
        RECT  0 0 168.7 99.12 ;
      LAYER via1 ;
        RECT  0 0 168.7 99.12 ;
      LAYER metal1 ;
        RECT  0 0 168.7 99.12 ;
    END
END fake_macro_newblue1_o330275

MACRO fake_macro_newblue1_o330276
    CLASS BLOCK ;
    SIZE 11.76 BY 252 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.765 9.555 128.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 123.165 10.115 123.235 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 118.965 10.115 119.035 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.725 9.555 130.795 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.965 1.155 224.035 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.925 1.155 176.995 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.645 1.155 239.715 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.125 1.155 216.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.085 1.155 169.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.245 1.155 161.315 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 158.445 9.555 158.515 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 134.645 10.115 134.715 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 138.565 10.115 138.635 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p249
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 252 ;
      LAYER metal2 ;
        RECT  0 0 11.76 252 ;
      LAYER via1 ;
        RECT  0 0 11.76 252 ;
      LAYER metal1 ;
        RECT  0 0 11.76 252 ;
    END
END fake_macro_newblue1_o330276

MACRO fake_macro_newblue1_o330277
    CLASS BLOCK ;
    SIZE 11.76 BY 252 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.765 9.555 128.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 123.165 10.115 123.235 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 118.965 10.115 119.035 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.725 9.555 130.795 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.925 1.155 176.995 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.245 1.155 161.315 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.085 1.155 169.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 158.445 9.555 158.515 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.125 1.155 216.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.645 1.155 239.715 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.965 1.155 224.035 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 134.645 10.115 134.715 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 138.565 10.115 138.635 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p249
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 252 ;
      LAYER metal2 ;
        RECT  0 0 11.76 252 ;
      LAYER via1 ;
        RECT  0 0 11.76 252 ;
      LAYER metal1 ;
        RECT  0 0 11.76 252 ;
    END
END fake_macro_newblue1_o330277

MACRO fake_macro_newblue1_o330278
    CLASS BLOCK ;
    SIZE 11.76 BY 252 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.725 9.555 130.795 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.765 9.555 128.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 123.165 10.115 123.235 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 118.965 10.115 119.035 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 158.445 9.555 158.515 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.645 1.155 239.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.925 1.155 176.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.965 1.155 224.035 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.125 1.155 216.195 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.245 1.155 161.315 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.085 1.155 169.155 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 134.645 10.115 134.715 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 138.565 10.115 138.635 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p249
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 252 ;
      LAYER metal2 ;
        RECT  0 0 11.76 252 ;
      LAYER via1 ;
        RECT  0 0 11.76 252 ;
      LAYER metal1 ;
        RECT  0 0 11.76 252 ;
    END
END fake_macro_newblue1_o330278

MACRO fake_macro_newblue1_o330279
    CLASS BLOCK ;
    SIZE 11.76 BY 252 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.725 9.555 130.795 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.765 9.555 128.835 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 123.165 10.115 123.235 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 118.965 10.115 119.035 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 158.445 9.555 158.515 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.085 1.155 169.155 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.245 1.155 161.315 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.925 1.155 176.995 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.125 1.155 216.195 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.645 1.155 239.715 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.965 1.155 224.035 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 134.645 10.115 134.715 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 138.565 10.115 138.635 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p249
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 252 ;
      LAYER metal2 ;
        RECT  0 0 11.76 252 ;
      LAYER via1 ;
        RECT  0 0 11.76 252 ;
      LAYER metal1 ;
        RECT  0 0 11.76 252 ;
    END
END fake_macro_newblue1_o330279

MACRO fake_macro_newblue1_o330280
    CLASS BLOCK ;
    SIZE 15.68 BY 142.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.885 13.475 73.955 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 68.285 14.035 68.355 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 64.085 14.035 64.155 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 71.365 1.155 71.435 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.245 1.155 70.315 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.845 13.475 75.915 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.565 13.475 75.635 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.285 1.155 110.355 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.645 1.155 127.715 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.845 1.155 82.915 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.805 1.155 21.875 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.765 1.155 79.835 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.685 1.155 83.755 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 103.565 13.475 103.635 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p75
    PIN p76
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p77
    PIN p78
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p79
    PIN p80
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p81
    PIN p82
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 79.765 14.035 79.835 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 83.685 14.035 83.755 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.325 1.155 80.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.245 1.155 84.315 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p139
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER via1 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal1 ;
        RECT  0 0 15.68 142.8 ;
    END
END fake_macro_newblue1_o330280

MACRO fake_macro_newblue1_o330281
    CLASS BLOCK ;
    SIZE 15.68 BY 142.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.845 13.475 75.915 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.885 13.475 73.955 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 68.285 14.035 68.355 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 64.085 14.035 64.155 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 71.365 1.155 71.435 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.245 1.155 70.315 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 103.565 13.475 103.635 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.565 13.475 75.635 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.805 1.155 21.875 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.845 1.155 82.915 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.645 1.155 127.715 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.285 1.155 110.355 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.765 1.155 79.835 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.685 1.155 83.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 79.765 14.035 79.835 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 83.685 14.035 83.755 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.325 1.155 80.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.245 1.155 84.315 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p139
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER via1 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal1 ;
        RECT  0 0 15.68 142.8 ;
    END
END fake_macro_newblue1_o330281

MACRO fake_macro_newblue1_o330282
    CLASS BLOCK ;
    SIZE 168.56 BY 99.12 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  165.165 97.125 165.235 97.195 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.005 97.125 159.075 97.195 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  156.205 97.125 156.275 97.195 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  154.525 97.125 154.595 97.195 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.845 97.125 152.915 97.195 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.165 97.125 151.235 97.195 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.925 97.125 148.995 97.195 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.245 97.125 147.315 97.195 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.565 97.125 145.635 97.195 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  143.885 97.125 143.955 97.195 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.725 97.125 137.795 97.195 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 97.125 136.115 97.195 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.805 97.125 133.875 97.195 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.125 97.125 132.195 97.195 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  130.445 97.125 130.515 97.195 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  128.765 97.125 128.835 97.195 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  126.525 97.125 126.595 97.195 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  124.845 97.125 124.915 97.195 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 97.125 122.115 97.195 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 97.125 120.435 97.195 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.685 97.125 118.755 97.195 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 97.125 117.075 97.195 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.765 97.125 114.835 97.195 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.085 97.125 113.155 97.195 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  111.405 97.125 111.475 97.195 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  109.725 97.125 109.795 97.195 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.565 97.125 103.635 97.195 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.885 97.125 101.955 97.195 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.645 97.125 99.715 97.195 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.965 97.125 98.035 97.195 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 97.125 96.355 97.195 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 97.125 94.675 97.195 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  92.365 97.125 92.435 97.195 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 97.125 90.755 97.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.885 97.125 87.955 97.195 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 97.125 86.275 97.195 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  84.525 97.125 84.595 97.195 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 97.125 82.915 97.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 97.125 80.675 97.195 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 97.125 78.995 97.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.245 97.125 77.315 97.195 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 97.125 75.635 97.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 97.125 69.475 97.195 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 97.125 67.795 97.195 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 97.125 65.555 97.195 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 97.125 63.875 97.195 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.125 97.125 62.195 97.195 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 97.125 60.515 97.195 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 97.125 58.275 97.195 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 97.125 56.595 97.195 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.725 97.125 53.795 97.195 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 97.125 52.115 97.195 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 97.125 50.435 97.195 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 97.125 48.755 97.195 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  46.445 97.125 46.515 97.195 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 97.125 44.835 97.195 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 97.125 43.155 97.195 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 97.125 41.475 97.195 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 97.125 35.315 97.195 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 97.125 33.635 97.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.325 97.125 31.395 97.195 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 97.125 29.715 97.195 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 97.125 28.035 97.195 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 97.125 26.355 97.195 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.045 97.125 24.115 97.195 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 97.125 22.435 97.195 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 93.205 12.355 93.275 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 96.845 6.755 96.915 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 93.205 16.275 93.275 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.085 93.205 15.155 93.275 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 98.805 12.355 98.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 86.765 3.395 86.835 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 92.085 5.635 92.155 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 85.645 2.275 85.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 93.205 14.595 93.275 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 76.405 3.955 76.475 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 78.645 3.395 78.715 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 78.645 3.955 78.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 80.885 3.395 80.955 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 80.885 3.955 80.955 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 67.445 3.395 67.515 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 67.445 3.955 67.515 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 69.685 3.395 69.755 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 69.685 3.955 69.755 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 71.925 3.395 71.995 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 71.925 3.955 71.995 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 74.165 3.395 74.235 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 74.165 3.955 74.235 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 76.405 3.395 76.475 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 98.805 3.955 98.875 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 78.925 4.515 78.995 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 67.725 4.515 67.795 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 67.165 4.515 67.235 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 69.965 4.515 70.035 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 69.405 4.515 69.475 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 72.205 4.515 72.275 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 71.645 4.515 71.715 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 85.925 12.915 85.995 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 97.125 22.995 97.195 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 97.125 25.235 97.195 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 97.125 26.915 97.195 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 97.125 28.595 97.195 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 97.125 30.275 97.195 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 97.125 32.515 97.195 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 97.125 34.195 97.195 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 97.125 35.875 97.195 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 97.125 42.035 97.195 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 97.125 43.715 97.195 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 97.125 45.395 97.195 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 97.125 47.635 97.195 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 97.125 49.315 97.195 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 97.125 50.995 97.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 97.125 52.675 97.195 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 97.125 54.915 97.195 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 97.125 57.155 97.195 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 97.125 59.395 97.195 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 97.125 61.075 97.195 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 97.125 62.755 97.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 97.125 64.435 97.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 97.125 66.675 97.195 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 97.125 68.355 97.195 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 97.125 70.035 97.195 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 97.125 76.195 97.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 97.125 77.875 97.195 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 97.125 79.555 97.195 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 97.125 81.795 97.195 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 97.125 83.475 97.195 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 97.125 85.155 97.195 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 97.125 86.835 97.195 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 97.125 89.075 97.195 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 97.125 91.315 97.195 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 97.125 93.555 97.195 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 97.125 95.235 97.195 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 97.125 96.915 97.195 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 97.125 98.595 97.195 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 97.125 100.835 97.195 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 97.125 102.515 97.195 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.125 97.125 104.195 97.195 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.285 97.125 110.355 97.195 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  111.965 97.125 112.035 97.195 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.645 97.125 113.715 97.195 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  115.885 97.125 115.955 97.195 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.565 97.125 117.635 97.195 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.245 97.125 119.315 97.195 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 97.125 120.995 97.195 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  123.165 97.125 123.235 97.195 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.405 97.125 125.475 97.195 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  127.645 97.125 127.715 97.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.325 97.125 129.395 97.195 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  131.005 97.125 131.075 97.195 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.685 97.125 132.755 97.195 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.925 97.125 134.995 97.195 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.605 97.125 136.675 97.195 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  138.285 97.125 138.355 97.195 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  144.445 97.125 144.515 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  146.125 97.125 146.195 97.195 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.805 97.125 147.875 97.195 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  150.045 97.125 150.115 97.195 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.725 97.125 151.795 97.195 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  153.405 97.125 153.475 97.195 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.085 97.125 155.155 97.195 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  157.325 97.125 157.395 97.195 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 97.125 159.635 97.195 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  165.725 97.125 165.795 97.195 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 96.845 11.795 96.915 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 92.365 7.875 92.435 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 86.765 3.955 86.835 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 85.365 2.275 85.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 80.605 23.555 80.675 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 80.605 25.235 80.675 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 80.605 27.475 80.675 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 80.605 29.155 80.675 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 80.605 30.835 80.675 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 80.605 32.515 80.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 80.605 34.755 80.675 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 80.605 36.435 80.675 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 80.605 42.595 80.675 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 80.605 44.275 80.675 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 80.605 45.955 80.675 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 80.605 47.635 80.675 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 80.605 49.875 80.675 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 80.605 51.555 80.675 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 80.605 53.235 80.675 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 80.605 54.915 80.675 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 80.605 57.715 80.675 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 80.605 59.395 80.675 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 80.605 61.635 80.675 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.245 80.605 63.315 80.675 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 80.605 64.995 80.675 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 80.605 66.675 80.675 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 80.605 68.915 80.675 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 80.605 70.595 80.675 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 80.605 76.755 80.675 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.365 80.605 78.435 80.675 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 80.605 80.115 80.675 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 80.605 81.795 80.675 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 80.605 84.035 80.675 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.645 80.605 85.715 80.675 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 80.605 87.395 80.675 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 80.605 89.075 80.675 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 80.605 91.875 80.675 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 80.605 93.555 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 80.605 95.795 80.675 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 80.605 97.475 80.675 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 80.605 99.155 80.675 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 80.605 100.835 80.675 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 80.605 103.075 80.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.685 80.605 104.755 80.675 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.845 80.605 110.915 80.675 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  112.525 80.605 112.595 80.675 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.205 80.605 114.275 80.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  115.885 80.605 115.955 80.675 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.125 80.605 118.195 80.675 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 80.605 119.875 80.675 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 80.605 121.555 80.675 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  123.165 80.605 123.235 80.675 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 80.605 126.035 80.675 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  127.645 80.605 127.715 80.675 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.885 80.605 129.955 80.675 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  131.565 80.605 131.635 80.675 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 80.605 133.315 80.675 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.925 80.605 134.995 80.675 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.165 80.605 137.235 80.675 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  138.845 80.605 138.915 80.675 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.005 80.605 145.075 80.675 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  146.685 80.605 146.755 80.675 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.365 80.605 148.435 80.675 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  150.045 80.605 150.115 80.675 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.285 80.605 152.355 80.675 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  153.965 80.605 154.035 80.675 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.645 80.605 155.715 80.675 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  157.325 80.605 157.395 80.675 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.125 80.605 160.195 80.675 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  166.285 80.605 166.355 80.675 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 98.805 2.275 98.875 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 78.645 10.675 78.715 ;
        END
    END p235
    OBS
      LAYER via2 ;
        RECT  0 0 168.7 99.12 ;
      LAYER metal2 ;
        RECT  0 0 168.7 99.12 ;
      LAYER via1 ;
        RECT  0 0 168.7 99.12 ;
      LAYER metal1 ;
        RECT  0 0 168.7 99.12 ;
    END
END fake_macro_newblue1_o330282

MACRO fake_macro_newblue1_o330283
    CLASS BLOCK ;
    SIZE 168.56 BY 99.12 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 93.205 12.355 93.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 96.845 6.755 96.915 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 93.205 16.275 93.275 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.085 93.205 15.155 93.275 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 98.805 12.355 98.875 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 86.765 3.395 86.835 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 85.645 2.275 85.715 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 93.205 14.595 93.275 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 76.405 3.955 76.475 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 78.645 3.395 78.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 78.645 3.955 78.715 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 80.885 3.395 80.955 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 80.885 3.955 80.955 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 67.445 3.395 67.515 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 67.445 3.955 67.515 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 69.685 3.395 69.755 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 69.685 3.955 69.755 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 71.925 3.395 71.995 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 71.925 3.955 71.995 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 74.165 3.395 74.235 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 74.165 3.955 74.235 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 76.405 3.395 76.475 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 96.845 11.795 96.915 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 92.365 7.875 92.435 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 98.805 3.955 98.875 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 78.925 4.515 78.995 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 67.725 4.515 67.795 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 67.165 4.515 67.235 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 69.965 4.515 70.035 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 69.405 4.515 69.475 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 72.205 4.515 72.275 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  4.445 71.645 4.515 71.715 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  109.725 97.125 109.795 97.195 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 97.125 96.355 97.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 97.125 86.275 97.195 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.245 97.125 77.315 97.195 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 97.125 63.875 97.195 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.725 97.125 53.795 97.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 97.125 44.835 97.195 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.325 97.125 31.395 97.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 97.125 22.435 97.195 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.845 97.125 152.915 97.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  143.885 97.125 143.955 97.195 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  130.445 97.125 130.515 97.195 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 97.125 120.435 97.195 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  111.405 97.125 111.475 97.195 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.965 97.125 98.035 97.195 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.885 97.125 87.955 97.195 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 97.125 78.995 97.195 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 97.125 65.555 97.195 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 97.125 56.595 97.195 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  46.445 97.125 46.515 97.195 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 97.125 33.635 97.195 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.045 97.125 24.115 97.195 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.005 97.125 159.075 97.195 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  156.205 97.125 156.275 97.195 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  154.525 97.125 154.595 97.195 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.925 97.125 148.995 97.195 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.565 97.125 145.635 97.195 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.725 97.125 137.795 97.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 97.125 136.115 97.195 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.125 97.125 132.195 97.195 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 97.125 122.115 97.195 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 97.125 117.075 97.195 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.765 97.125 114.835 97.195 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.885 97.125 101.955 97.195 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  92.365 97.125 92.435 97.195 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 97.125 69.475 97.195 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 97.125 60.515 97.195 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 97.125 52.115 97.195 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 97.125 26.355 97.195 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.245 97.125 147.315 97.195 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.805 97.125 133.875 97.195 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.565 97.125 103.635 97.195 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  84.525 97.125 84.595 97.195 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 97.125 67.795 97.195 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 97.125 48.755 97.195 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 97.125 41.475 97.195 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 97.125 29.715 97.195 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 97.125 28.035 97.195 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.165 97.125 151.235 97.195 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  128.765 97.125 128.835 97.195 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  126.525 97.125 126.595 97.195 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  124.845 97.125 124.915 97.195 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.685 97.125 118.755 97.195 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.645 97.125 99.715 97.195 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 97.125 94.675 97.195 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 97.125 90.755 97.195 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 97.125 82.915 97.195 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 97.125 80.675 97.195 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 97.125 75.635 97.195 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.125 97.125 62.195 97.195 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 97.125 58.275 97.195 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 97.125 50.435 97.195 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 97.125 43.155 97.195 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 97.125 35.315 97.195 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  165.165 97.125 165.235 97.195 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.085 97.125 113.155 97.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 85.925 12.915 85.995 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 97.125 22.995 97.195 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 97.125 25.235 97.195 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 97.125 26.915 97.195 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 97.125 28.595 97.195 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 97.125 30.275 97.195 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 97.125 32.515 97.195 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 97.125 34.195 97.195 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 97.125 35.875 97.195 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 97.125 42.035 97.195 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 97.125 43.715 97.195 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 97.125 45.395 97.195 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 97.125 47.635 97.195 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 97.125 49.315 97.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 97.125 50.995 97.195 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 97.125 52.675 97.195 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 97.125 54.915 97.195 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 97.125 57.155 97.195 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 97.125 59.395 97.195 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 97.125 61.075 97.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 97.125 62.755 97.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 97.125 64.435 97.195 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 97.125 66.675 97.195 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 97.125 68.355 97.195 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 97.125 70.035 97.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 97.125 76.195 97.195 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 97.125 77.875 97.195 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 97.125 79.555 97.195 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 97.125 81.795 97.195 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 97.125 83.475 97.195 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 97.125 85.155 97.195 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 97.125 86.835 97.195 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 97.125 89.075 97.195 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 97.125 91.315 97.195 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 97.125 93.555 97.195 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 97.125 95.235 97.195 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 97.125 96.915 97.195 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 97.125 98.595 97.195 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 97.125 100.835 97.195 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 97.125 102.515 97.195 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.125 97.125 104.195 97.195 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.285 97.125 110.355 97.195 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  111.965 97.125 112.035 97.195 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.645 97.125 113.715 97.195 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  115.885 97.125 115.955 97.195 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.565 97.125 117.635 97.195 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.245 97.125 119.315 97.195 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 97.125 120.995 97.195 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  123.165 97.125 123.235 97.195 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.405 97.125 125.475 97.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  127.645 97.125 127.715 97.195 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.325 97.125 129.395 97.195 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  131.005 97.125 131.075 97.195 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.685 97.125 132.755 97.195 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.925 97.125 134.995 97.195 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.605 97.125 136.675 97.195 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  138.285 97.125 138.355 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  144.445 97.125 144.515 97.195 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  146.125 97.125 146.195 97.195 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.805 97.125 147.875 97.195 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  150.045 97.125 150.115 97.195 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.725 97.125 151.795 97.195 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  153.405 97.125 153.475 97.195 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.085 97.125 155.155 97.195 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  157.325 97.125 157.395 97.195 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 97.125 159.635 97.195 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  165.725 97.125 165.795 97.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 92.085 5.635 92.155 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 86.765 3.955 86.835 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 85.365 2.275 85.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 80.605 23.555 80.675 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 80.605 25.235 80.675 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 80.605 27.475 80.675 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 80.605 29.155 80.675 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 80.605 30.835 80.675 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  32.445 80.605 32.515 80.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 80.605 34.755 80.675 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.365 80.605 36.435 80.675 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 80.605 42.595 80.675 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 80.605 44.275 80.675 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 80.605 45.955 80.675 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 80.605 47.635 80.675 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 80.605 49.875 80.675 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 80.605 51.555 80.675 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 80.605 53.235 80.675 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.845 80.605 54.915 80.675 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 80.605 57.715 80.675 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 80.605 59.395 80.675 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 80.605 61.635 80.675 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.245 80.605 63.315 80.675 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 80.605 64.995 80.675 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 80.605 66.675 80.675 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 80.605 68.915 80.675 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 80.605 70.595 80.675 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 80.605 76.755 80.675 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.365 80.605 78.435 80.675 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 80.605 80.115 80.675 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 80.605 81.795 80.675 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 80.605 84.035 80.675 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.645 80.605 85.715 80.675 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 80.605 87.395 80.675 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 80.605 89.075 80.675 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 80.605 91.875 80.675 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 80.605 93.555 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 80.605 95.795 80.675 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 80.605 97.475 80.675 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 80.605 99.155 80.675 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 80.605 100.835 80.675 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 80.605 103.075 80.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.685 80.605 104.755 80.675 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.845 80.605 110.915 80.675 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  112.525 80.605 112.595 80.675 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.205 80.605 114.275 80.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  115.885 80.605 115.955 80.675 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.125 80.605 118.195 80.675 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 80.605 119.875 80.675 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 80.605 121.555 80.675 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  123.165 80.605 123.235 80.675 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 80.605 126.035 80.675 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  127.645 80.605 127.715 80.675 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.885 80.605 129.955 80.675 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  131.565 80.605 131.635 80.675 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 80.605 133.315 80.675 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.925 80.605 134.995 80.675 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.165 80.605 137.235 80.675 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  138.845 80.605 138.915 80.675 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.005 80.605 145.075 80.675 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  146.685 80.605 146.755 80.675 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.365 80.605 148.435 80.675 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  150.045 80.605 150.115 80.675 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.285 80.605 152.355 80.675 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  153.965 80.605 154.035 80.675 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.645 80.605 155.715 80.675 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  157.325 80.605 157.395 80.675 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.125 80.605 160.195 80.675 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  166.285 80.605 166.355 80.675 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 98.805 2.275 98.875 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 78.645 10.675 78.715 ;
        END
    END p235
    OBS
      LAYER via2 ;
        RECT  0 0 168.7 99.12 ;
      LAYER metal2 ;
        RECT  0 0 168.7 99.12 ;
      LAYER via1 ;
        RECT  0 0 168.7 99.12 ;
      LAYER metal1 ;
        RECT  0 0 168.7 99.12 ;
    END
END fake_macro_newblue1_o330283

MACRO fake_macro_newblue1_o330284
    CLASS BLOCK ;
    SIZE 11.76 BY 252 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.725 9.555 130.795 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.765 9.555 128.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 123.165 10.115 123.235 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 118.965 10.115 119.035 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 158.445 9.555 158.515 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.965 1.155 224.035 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.925 1.155 176.995 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.085 1.155 169.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.245 1.155 161.315 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.645 1.155 239.715 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.125 1.155 216.195 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 134.645 10.115 134.715 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 138.565 10.115 138.635 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p249
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 252 ;
      LAYER metal2 ;
        RECT  0 0 11.76 252 ;
      LAYER via1 ;
        RECT  0 0 11.76 252 ;
      LAYER metal1 ;
        RECT  0 0 11.76 252 ;
    END
END fake_macro_newblue1_o330284

MACRO fake_macro_newblue1_o330285
    CLASS BLOCK ;
    SIZE 11.76 BY 252 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.725 9.555 130.795 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.765 9.555 128.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 123.165 10.115 123.235 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 118.965 10.115 119.035 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 158.445 9.555 158.515 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.925 1.155 176.995 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.245 1.155 161.315 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.085 1.155 169.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.125 1.155 216.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.645 1.155 239.715 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.965 1.155 224.035 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 134.645 10.115 134.715 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 138.565 10.115 138.635 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p249
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 252 ;
      LAYER metal2 ;
        RECT  0 0 11.76 252 ;
      LAYER via1 ;
        RECT  0 0 11.76 252 ;
      LAYER metal1 ;
        RECT  0 0 11.76 252 ;
    END
END fake_macro_newblue1_o330285

MACRO fake_macro_newblue1_o330286
    CLASS BLOCK ;
    SIZE 11.76 BY 252 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.725 9.555 130.795 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.765 9.555 128.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 123.165 10.115 123.235 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 118.965 10.115 119.035 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 158.445 9.555 158.515 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.645 1.155 239.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.925 1.155 176.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.965 1.155 224.035 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.125 1.155 216.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.245 1.155 161.315 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.085 1.155 169.155 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 134.645 10.115 134.715 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 138.565 10.115 138.635 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p249
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 252 ;
      LAYER metal2 ;
        RECT  0 0 11.76 252 ;
      LAYER via1 ;
        RECT  0 0 11.76 252 ;
      LAYER metal1 ;
        RECT  0 0 11.76 252 ;
    END
END fake_macro_newblue1_o330286

MACRO fake_macro_newblue1_o330287
    CLASS BLOCK ;
    SIZE 11.76 BY 252 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.725 9.555 130.795 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.765 9.555 128.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 123.165 10.115 123.235 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 118.965 10.115 119.035 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 158.445 9.555 158.515 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.085 1.155 169.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.245 1.155 161.315 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.925 1.155 176.995 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.125 1.155 216.195 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.645 1.155 239.715 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.965 1.155 224.035 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 134.645 10.115 134.715 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 138.565 10.115 138.635 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p249
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 252 ;
      LAYER metal2 ;
        RECT  0 0 11.76 252 ;
      LAYER via1 ;
        RECT  0 0 11.76 252 ;
      LAYER metal1 ;
        RECT  0 0 11.76 252 ;
    END
END fake_macro_newblue1_o330287

MACRO fake_macro_newblue1_o330288
    CLASS BLOCK ;
    SIZE 15.68 BY 142.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.845 13.475 75.915 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.885 13.475 73.955 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 68.285 14.035 68.355 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 64.085 14.035 64.155 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 71.365 1.155 71.435 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.245 1.155 70.315 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 103.565 13.475 103.635 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.565 13.475 75.635 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.285 1.155 110.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.645 1.155 127.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.845 1.155 82.915 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.805 1.155 21.875 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.765 1.155 79.835 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.685 1.155 83.755 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p75
    PIN p76
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p77
    PIN p78
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p79
    PIN p80
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p81
    PIN p82
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 79.765 14.035 79.835 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 83.685 14.035 83.755 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.325 1.155 80.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.245 1.155 84.315 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p139
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER via1 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal1 ;
        RECT  0 0 15.68 142.8 ;
    END
END fake_macro_newblue1_o330288

MACRO fake_macro_newblue1_o330289
    CLASS BLOCK ;
    SIZE 15.68 BY 142.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.845 13.475 75.915 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.885 13.475 73.955 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 68.285 14.035 68.355 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 64.085 14.035 64.155 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 71.365 1.155 71.435 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.245 1.155 70.315 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 103.565 13.475 103.635 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.565 13.475 75.635 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.805 1.155 21.875 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.845 1.155 82.915 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.645 1.155 127.715 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.285 1.155 110.355 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.765 1.155 79.835 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.685 1.155 83.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 79.765 14.035 79.835 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 83.685 14.035 83.755 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.325 1.155 80.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.245 1.155 84.315 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p139
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER via1 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal1 ;
        RECT  0 0 15.68 142.8 ;
    END
END fake_macro_newblue1_o330289

MACRO fake_macro_newblue1_o330290
    CLASS BLOCK ;
    SIZE 55.44 BY 31.92 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 29.365 13.475 29.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 28.245 1.715 28.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.365 6.755 29.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 29.365 11.235 29.435 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 29.365 15.715 29.435 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 31.605 15.715 31.675 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 29.365 10.675 29.435 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 29.365 6.195 29.435 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 27.405 1.715 27.475 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 24.885 1.715 24.955 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 31.605 6.755 31.675 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 31.605 11.235 31.675 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 29.365 21.875 29.435 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 5.845 24.675 5.915 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 5.565 22.435 5.635 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 20.125 53.235 20.195 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 29.365 21.315 29.435 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.005 1.715 12.075 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 6.125 12.355 6.195 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 6.125 22.995 6.195 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 19.005 53.235 19.075 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 19.565 47.635 19.635 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  20.125 29.365 20.195 29.435 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 29.365 22.995 29.435 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 22.365 53.235 22.435 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 24.045 53.235 24.115 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 25.725 53.235 25.795 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 27.405 53.235 27.475 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 29.085 53.235 29.155 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 3.885 53.235 3.955 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 5.565 53.235 5.635 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 7.245 53.235 7.315 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 8.925 53.235 8.995 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 10.605 53.235 10.675 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 12.285 53.235 12.355 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 13.965 53.235 14.035 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 15.645 53.235 15.715 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 17.325 53.235 17.395 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 24.045 1.715 24.115 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  20.125 31.605 20.195 31.675 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 20.125 48.755 20.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.605 31.605 10.675 31.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 29.085 15.715 29.155 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 29.365 14.035 29.435 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 20.685 49.315 20.755 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 21.245 53.235 21.315 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 29.645 16.275 29.715 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 29.365 45.395 29.435 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 29.365 45.955 29.435 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.165 29.365 25.235 29.435 ;
        END
    END p50
    OBS
      LAYER via2 ;
        RECT  0 0 55.44 31.92 ;
      LAYER metal2 ;
        RECT  0 0 55.44 31.92 ;
      LAYER via1 ;
        RECT  0 0 55.44 31.92 ;
      LAYER metal1 ;
        RECT  0 0 55.44 31.92 ;
    END
END fake_macro_newblue1_o330290

MACRO fake_macro_newblue1_o330327
    CLASS BLOCK ;
    SIZE 122.92 BY 189.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.885 1.155 3.955 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.365 1.155 8.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.685 1.155 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.845 1.155 12.915 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.525 1.155 14.595 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.325 1.155 17.395 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.645 1.155 15.715 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.805 1.155 21.875 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 20.125 1.155 20.195 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.285 1.155 26.355 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 24.605 1.155 24.675 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.765 1.155 30.835 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.085 1.155 29.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.245 1.155 35.315 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 36.925 1.155 36.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.725 1.155 39.795 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.045 1.155 38.115 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 44.205 1.155 44.275 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.525 1.155 42.595 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 48.685 1.155 48.755 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.365 1.155 50.435 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.485 1.155 51.555 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.645 1.155 57.715 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.325 1.155 59.395 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.125 1.155 62.195 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 60.445 1.155 60.515 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.605 1.155 66.675 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 71.085 1.155 71.155 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.405 1.155 69.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 75.565 1.155 75.635 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.885 1.155 73.955 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.045 1.155 80.115 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.365 1.155 78.435 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 114.485 1.155 114.555 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.125 1.155 125.195 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.605 1.155 129.675 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.405 1.155 132.475 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.085 1.155 134.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 143.045 3.395 143.115 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.845 1.155 145.915 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.525 1.155 147.595 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 152.005 1.155 152.075 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 156.485 1.155 156.555 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.285 1.155 159.355 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 163.765 1.155 163.835 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 165.445 1.155 165.515 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.245 1.155 168.315 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 172.725 1.155 172.795 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.205 1.155 177.275 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.885 1.155 178.955 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 183.365 1.155 183.435 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 187.845 1.155 187.915 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.245 84.525 119.315 84.595 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 85.645 120.435 85.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.245 88.725 119.315 88.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.405 1.155 97.475 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.405 1.155 83.475 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 94.885 2.275 94.955 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 101.045 119.875 101.115 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 105.525 120.995 105.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.685 1.155 83.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 94.885 2.835 94.955 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 101.325 119.875 101.395 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 105.805 120.995 105.875 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.765 1.155 86.835 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.685 1.155 90.755 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.645 1.155 99.715 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.925 1.155 106.995 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.885 1.155 87.955 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.405 1.155 118.475 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 98.245 1.155 98.315 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.685 1.155 104.755 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.965 1.155 98.035 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 89.565 1.715 89.635 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 98.245 1.715 98.315 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 104.685 1.715 104.755 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.245 112.245 119.315 112.315 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.205 1.155 184.275 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 187.005 2.835 187.075 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 179.725 1.155 179.795 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 182.525 2.835 182.595 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 178.045 1.715 178.115 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 178.045 2.835 178.115 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.765 1.155 170.835 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 173.565 2.835 173.635 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.285 1.155 166.355 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 169.085 2.835 169.155 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 161.805 1.155 161.875 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 164.605 2.835 164.675 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 157.325 1.155 157.395 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 160.125 2.835 160.195 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 155.645 1.715 155.715 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 155.645 2.835 155.715 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 148.365 1.155 148.435 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 151.165 2.835 151.235 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.885 1.155 143.955 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 146.685 2.835 146.755 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 142.205 1.715 142.275 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 142.205 2.835 142.275 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.925 1.155 134.995 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 137.725 2.835 137.795 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.445 1.155 130.515 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 133.245 2.835 133.315 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.965 1.155 126.035 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 128.765 2.835 128.835 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.485 1.155 121.555 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 124.285 2.835 124.355 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.005 1.155 117.075 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 119.805 2.835 119.875 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.525 1.155 112.595 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 115.325 2.835 115.395 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 110.845 2.835 110.915 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 82.285 1.715 82.355 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 82.285 2.835 82.355 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 77.805 1.715 77.875 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 77.805 2.835 77.875 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 73.325 1.715 73.395 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 73.325 2.835 73.395 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 68.845 1.715 68.915 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 68.845 2.835 68.915 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 64.365 1.715 64.435 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 64.365 2.835 64.435 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 59.885 1.715 59.955 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 59.885 2.835 59.955 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 55.405 1.715 55.475 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 55.405 2.835 55.475 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 50.925 1.715 50.995 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 50.925 2.835 50.995 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 46.445 1.715 46.515 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 46.445 2.835 46.515 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 41.965 1.715 42.035 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 41.965 2.835 42.035 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 37.485 1.715 37.555 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 37.485 2.835 37.555 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 33.005 1.715 33.075 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 33.005 2.835 33.075 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 28.525 1.715 28.595 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 28.525 2.835 28.595 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 24.045 1.715 24.115 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 24.045 2.835 24.115 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 19.565 1.715 19.635 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 19.565 2.835 19.635 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 15.085 1.715 15.155 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 15.085 2.835 15.155 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 10.605 1.715 10.675 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 10.605 2.835 10.675 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 6.125 1.715 6.195 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 6.125 2.835 6.195 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.245 85.365 119.315 85.435 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 97.965 1.715 98.035 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 187.565 120.995 187.635 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 189.525 120.995 189.595 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 183.085 120.995 183.155 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 183.365 121.555 183.435 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 177.205 120.995 177.275 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 178.605 120.995 178.675 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 174.125 120.995 174.195 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 174.405 121.555 174.475 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 169.645 120.995 169.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 169.925 121.555 169.995 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 165.165 120.995 165.235 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 165.445 121.555 165.515 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 160.685 120.995 160.755 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 160.965 121.555 161.035 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 156.205 120.995 156.275 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 156.485 121.555 156.555 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 151.725 120.995 151.795 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 152.005 121.555 152.075 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 147.245 120.995 147.315 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 147.525 121.555 147.595 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 141.365 120.995 141.435 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 141.925 120.995 141.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 138.285 120.995 138.355 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 138.565 121.555 138.635 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 133.805 120.995 133.875 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 134.085 121.555 134.155 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 129.325 120.995 129.395 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 129.605 121.555 129.675 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 124.845 120.995 124.915 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 125.125 121.555 125.195 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 120.365 120.995 120.435 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 120.645 121.555 120.715 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 115.885 120.995 115.955 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 116.165 121.555 116.235 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 111.405 120.995 111.475 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 111.685 121.555 111.755 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 81.445 120.995 81.515 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 83.405 120.995 83.475 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 76.965 120.995 77.035 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 77.245 121.555 77.315 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 72.485 120.995 72.555 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 72.765 121.555 72.835 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 68.005 120.995 68.075 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 68.285 121.555 68.355 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 63.525 120.995 63.595 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 63.805 121.555 63.875 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 59.045 120.995 59.115 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 59.325 121.555 59.395 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 54.565 120.995 54.635 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 54.845 121.555 54.915 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 50.085 120.995 50.155 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 50.365 121.555 50.435 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 45.605 120.995 45.675 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 45.885 121.555 45.955 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 41.125 120.995 41.195 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 41.405 121.555 41.475 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 36.645 120.995 36.715 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 34.685 120.995 34.755 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 32.165 120.995 32.235 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 32.445 121.555 32.515 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 27.685 120.995 27.755 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 27.965 121.555 28.035 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 23.205 120.995 23.275 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 23.485 121.555 23.555 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 18.725 120.995 18.795 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 19.005 121.555 19.075 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 14.245 120.995 14.315 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 14.525 121.555 14.595 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 9.765 120.995 9.835 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 10.045 121.555 10.115 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 5.285 120.995 5.355 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 5.565 121.555 5.635 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.725 1.155 186.795 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.285 1.155 173.355 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 164.325 1.155 164.395 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.845 1.155 159.915 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.365 1.155 155.435 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 169.925 1.715 169.995 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.445 1.155 137.515 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.965 1.155 133.035 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.485 1.155 128.555 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.565 1.155 110.635 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.485 1.155 79.555 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 75.005 1.155 75.075 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.525 1.155 70.595 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.045 1.155 66.115 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.565 1.155 61.635 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 52.605 1.155 52.675 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 48.125 1.155 48.195 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.645 1.155 43.715 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.165 1.155 39.235 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.685 1.155 34.755 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.205 1.155 30.275 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.725 1.155 25.795 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.245 1.155 21.315 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 16.765 1.155 16.835 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.285 1.155 12.355 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.805 1.155 7.875 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.325 1.155 3.395 ;
        END
    END p284
    OBS
      LAYER via2 ;
        RECT  0 0 122.92 189.84 ;
      LAYER metal2 ;
        RECT  0 0 122.92 189.84 ;
      LAYER via1 ;
        RECT  0 0 122.92 189.84 ;
      LAYER metal1 ;
        RECT  0 0 122.92 189.84 ;
    END
END fake_macro_newblue1_o330327

MACRO fake_macro_newblue1_o330440
    CLASS BLOCK ;
    SIZE 20.16 BY 273.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.765 143.605 16.835 143.675 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.525 1.155 147.595 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.445 1.155 151.515 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.365 1.155 155.435 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.285 1.155 159.355 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 163.205 1.155 163.275 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 167.125 1.155 167.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.045 1.155 171.115 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.965 1.155 175.035 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.885 1.155 178.955 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.805 1.155 182.875 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.725 1.155 186.795 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.645 1.155 190.715 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.565 1.155 194.635 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.485 1.155 198.555 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.405 1.155 202.475 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.325 1.155 206.395 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 210.245 1.155 210.315 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 214.165 1.155 214.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 218.085 1.155 218.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 222.005 1.155 222.075 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.925 1.155 225.995 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.845 1.155 229.915 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.765 1.155 233.835 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.685 1.155 237.755 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.605 1.155 241.675 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.525 1.155 245.595 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 249.445 1.155 249.515 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.365 1.155 253.435 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.285 1.155 257.355 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 261.205 1.155 261.275 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 265.125 1.155 265.195 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 269.045 1.155 269.115 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.525 1.155 35.595 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 98.245 1.155 98.315 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.765 1.155 121.835 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.685 1.155 125.755 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 148.365 1.155 148.435 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 152.285 1.155 152.355 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 156.205 1.155 156.275 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.125 1.155 160.195 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.365 1.155 162.435 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 167.965 1.155 168.035 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.885 1.155 171.955 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 175.805 1.155 175.875 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.045 1.155 178.115 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 183.645 1.155 183.715 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 187.565 1.155 187.635 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 191.485 1.155 191.555 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 195.405 1.155 195.475 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 199.325 1.155 199.395 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 203.245 1.155 203.315 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 207.165 1.155 207.235 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 211.085 1.155 211.155 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.325 1.155 213.395 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 218.925 1.155 218.995 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 222.845 1.155 222.915 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 226.765 1.155 226.835 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 230.685 1.155 230.755 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 234.605 1.155 234.675 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 238.525 1.155 238.595 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 242.445 1.155 242.515 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 246.365 1.155 246.435 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 250.285 1.155 250.355 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 254.205 1.155 254.275 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 258.125 1.155 258.195 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.285 1.155 264.355 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 269.885 1.155 269.955 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 144.725 1.155 144.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.765 171.325 16.835 171.395 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 142.765 17.955 142.835 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 141.645 17.955 141.715 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 136.885 17.955 136.955 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.085 1.155 127.155 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 141.365 1.155 141.435 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.045 1.155 136.115 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 126.805 17.955 126.875 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 140.805 1.155 140.875 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.485 1.155 135.555 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 154.525 17.955 154.595 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 144.445 1.155 144.515 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.685 1.155 132.755 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.605 1.155 129.675 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.045 1.155 262.115 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 3.045 17.955 3.115 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 2.765 18.515 2.835 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 6.965 17.955 7.035 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 6.405 18.515 6.475 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 10.885 17.955 10.955 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 10.605 18.515 10.675 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 14.805 17.955 14.875 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 14.245 18.515 14.315 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 18.725 17.955 18.795 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 18.165 18.515 18.235 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 22.645 17.955 22.715 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 22.365 18.515 22.435 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 25.445 17.955 25.515 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 26.285 18.515 26.355 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 30.485 17.955 30.555 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 29.925 18.515 29.995 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 33.285 17.955 33.355 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 34.125 18.515 34.195 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 38.325 17.955 38.395 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 37.765 18.515 37.835 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 42.245 17.955 42.315 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 41.685 18.515 41.755 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 46.165 17.955 46.235 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 45.885 18.515 45.955 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 50.085 17.955 50.155 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 49.525 18.515 49.595 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 54.005 17.955 54.075 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 53.445 18.515 53.515 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 57.925 17.955 57.995 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 57.645 18.515 57.715 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 61.845 17.955 61.915 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 61.565 18.515 61.635 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 65.765 17.955 65.835 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 65.205 18.515 65.275 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 69.685 17.955 69.755 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 69.405 18.515 69.475 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 73.605 17.955 73.675 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 73.325 18.515 73.395 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 76.405 17.955 76.475 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 77.245 18.515 77.315 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 81.445 17.955 81.515 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 81.165 18.515 81.235 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 84.245 17.955 84.315 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 84.805 18.515 84.875 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 89.285 17.955 89.355 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 88.725 18.515 88.795 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 93.205 17.955 93.275 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 92.925 18.515 92.995 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 97.125 17.955 97.195 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 96.845 18.515 96.915 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 101.045 17.955 101.115 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 100.485 18.515 100.555 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 104.965 17.955 105.035 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 104.685 18.515 104.755 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 108.885 17.955 108.955 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 108.325 18.515 108.395 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 112.805 17.955 112.875 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 112.525 18.515 112.595 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 116.725 17.955 116.795 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 116.445 18.515 116.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 119.525 17.955 119.595 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 120.365 18.515 120.435 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 124.565 17.955 124.635 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 124.285 18.515 124.355 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 147.805 17.955 147.875 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 146.685 18.515 146.755 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 151.725 17.955 151.795 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 150.605 18.515 150.675 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 155.645 17.955 155.715 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 154.525 18.515 154.595 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 159.565 17.955 159.635 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 158.445 18.515 158.515 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 163.485 17.955 163.555 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 162.365 18.515 162.435 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 167.405 17.955 167.475 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 166.285 18.515 166.355 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 171.045 17.955 171.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 170.205 18.515 170.275 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 175.245 17.955 175.315 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 174.125 18.515 174.195 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 178.885 17.955 178.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 179.445 18.515 179.515 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 183.085 17.955 183.155 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 181.965 18.515 182.035 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 186.725 17.955 186.795 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 187.285 18.515 187.355 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 190.925 17.955 190.995 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 189.805 18.515 189.875 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 194.845 17.955 194.915 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 193.725 18.515 193.795 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 198.765 17.955 198.835 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 197.645 18.515 197.715 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 202.685 17.955 202.755 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 201.565 18.515 201.635 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 206.605 17.955 206.675 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 205.485 18.515 205.555 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 210.525 17.955 210.595 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 209.405 18.515 209.475 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 214.445 17.955 214.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 213.325 18.515 213.395 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 218.365 17.955 218.435 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 217.245 18.515 217.315 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 222.005 17.955 222.075 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 221.165 18.515 221.235 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 226.205 17.955 226.275 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 225.085 18.515 225.155 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 230.125 17.955 230.195 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 230.405 18.515 230.475 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 234.045 17.955 234.115 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 232.925 18.515 232.995 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 237.965 17.955 238.035 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 236.845 18.515 236.915 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 241.885 17.955 241.955 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 240.765 18.515 240.835 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 245.805 17.955 245.875 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 244.685 18.515 244.755 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 249.725 17.955 249.795 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 248.605 18.515 248.675 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 253.645 17.955 253.715 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 252.525 18.515 252.595 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 257.565 17.955 257.635 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 256.445 18.515 256.515 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 261.485 17.955 261.555 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 260.365 18.515 260.435 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 265.125 17.955 265.195 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 264.285 18.515 264.355 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 269.325 17.955 269.395 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 268.205 18.515 268.275 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p285
    PIN p286
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p287
    PIN p288
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p289
    PIN p290
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p291
    PIN p292
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p293
    PIN p294
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p295
    PIN p296
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 148.085 1.155 148.155 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 152.005 1.155 152.075 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.925 1.155 155.995 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.845 1.155 159.915 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 163.765 1.155 163.835 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 167.685 1.155 167.755 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.605 1.155 171.675 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 175.525 1.155 175.595 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 179.445 1.155 179.515 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 183.365 1.155 183.435 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 187.285 1.155 187.355 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 191.205 1.155 191.275 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 195.125 1.155 195.195 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 199.045 1.155 199.115 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.965 1.155 203.035 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.885 1.155 206.955 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 210.805 1.155 210.875 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 214.725 1.155 214.795 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 218.645 1.155 218.715 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 222.565 1.155 222.635 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 226.485 1.155 226.555 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 230.405 1.155 230.475 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 234.325 1.155 234.395 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 238.245 1.155 238.315 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 242.165 1.155 242.235 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 246.085 1.155 246.155 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 250.005 1.155 250.075 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.925 1.155 253.995 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.845 1.155 257.915 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 261.765 1.155 261.835 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 265.685 1.155 265.755 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 269.605 1.155 269.675 ;
        END
    END p335
    OBS
      LAYER via2 ;
        RECT  0 0 20.16 273.84 ;
      LAYER metal2 ;
        RECT  0 0 20.16 273.84 ;
      LAYER via1 ;
        RECT  0 0 20.16 273.84 ;
      LAYER metal1 ;
        RECT  0 0 20.16 273.84 ;
    END
END fake_macro_newblue1_o330440

MACRO fake_macro_newblue1_o330441
    CLASS BLOCK ;
    SIZE 11.76 BY 268.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.525 1.155 35.595 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.005 1.155 61.075 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.645 1.155 78.715 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 94.325 1.155 94.395 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.125 1.155 104.195 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.965 1.155 112.035 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.685 1.155 125.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.085 1.155 155.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.925 1.155 162.995 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.765 1.155 170.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.605 1.155 178.675 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.445 1.155 186.515 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 188.685 1.155 188.755 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.285 1.155 194.355 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 196.525 1.155 196.595 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.125 1.155 202.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 204.365 1.155 204.435 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.965 1.155 210.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.805 1.155 217.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.645 1.155 225.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.485 1.155 233.555 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.325 1.155 241.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.085 1.155 253.155 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.325 1.155 255.395 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.925 1.155 260.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 263.165 1.155 263.235 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 131.005 10.115 131.075 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 126.805 10.115 126.875 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 136.605 9.555 136.675 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.325 1.155 136.395 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.565 9.555 138.635 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.285 9.555 138.355 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.245 1.155 252.315 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.165 1.155 256.235 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.085 1.155 260.155 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.005 1.155 264.075 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 166.285 9.555 166.355 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 120.645 10.115 120.715 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 124.565 10.115 124.635 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 252.245 10.115 252.315 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 256.165 10.115 256.235 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 260.085 10.115 260.155 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 264.005 10.115 264.075 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.805 1.155 252.875 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.645 1.155 260.715 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p265
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER via1 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal1 ;
        RECT  0 0 11.76 268.8 ;
    END
END fake_macro_newblue1_o330441

MACRO fake_macro_newblue1_o330442
    CLASS BLOCK ;
    SIZE 20.16 BY 273.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.765 143.605 16.835 143.675 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 142.765 17.955 142.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.965 1.155 175.035 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.805 1.155 182.875 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 210.245 1.155 210.315 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 218.085 1.155 218.155 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.925 1.155 225.995 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.685 1.155 237.755 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.365 1.155 253.435 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.285 1.155 257.355 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 261.205 1.155 261.275 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 265.125 1.155 265.195 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.525 1.155 35.595 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 98.245 1.155 98.315 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.765 1.155 121.835 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.685 1.155 125.755 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 148.365 1.155 148.435 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 152.285 1.155 152.355 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 156.205 1.155 156.275 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.125 1.155 160.195 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.365 1.155 162.435 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 167.965 1.155 168.035 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.885 1.155 171.955 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 175.805 1.155 175.875 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.045 1.155 178.115 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 183.645 1.155 183.715 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 187.565 1.155 187.635 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 191.485 1.155 191.555 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 195.405 1.155 195.475 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 199.325 1.155 199.395 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 203.245 1.155 203.315 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 207.165 1.155 207.235 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 211.085 1.155 211.155 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.325 1.155 213.395 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 218.925 1.155 218.995 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 222.845 1.155 222.915 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 226.765 1.155 226.835 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 230.685 1.155 230.755 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 234.605 1.155 234.675 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 238.525 1.155 238.595 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 242.445 1.155 242.515 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 246.365 1.155 246.435 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 250.285 1.155 250.355 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 254.205 1.155 254.275 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 258.125 1.155 258.195 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.045 1.155 262.115 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.285 1.155 264.355 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 269.885 1.155 269.955 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.085 1.155 127.155 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 126.805 17.955 126.875 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 154.525 17.955 154.595 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.605 1.155 129.675 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 144.725 1.155 144.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 141.645 17.955 141.715 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 136.885 17.955 136.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 141.365 1.155 141.435 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.045 1.155 136.115 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 140.805 1.155 140.875 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.485 1.155 135.555 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 144.445 1.155 144.515 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.685 1.155 132.755 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.765 171.325 16.835 171.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.525 1.155 147.595 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.445 1.155 151.515 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.365 1.155 155.435 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.285 1.155 159.355 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 163.205 1.155 163.275 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 167.125 1.155 167.195 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.045 1.155 171.115 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.885 1.155 178.955 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.725 1.155 186.795 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.645 1.155 190.715 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.565 1.155 194.635 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.485 1.155 198.555 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.405 1.155 202.475 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.325 1.155 206.395 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 214.165 1.155 214.235 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 222.005 1.155 222.075 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.845 1.155 229.915 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.765 1.155 233.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.605 1.155 241.675 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.525 1.155 245.595 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 249.445 1.155 249.515 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 269.045 1.155 269.115 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 3.045 17.955 3.115 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 2.765 18.515 2.835 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 6.965 17.955 7.035 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 6.405 18.515 6.475 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 10.885 17.955 10.955 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 10.605 18.515 10.675 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 14.805 17.955 14.875 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 14.245 18.515 14.315 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 18.725 17.955 18.795 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 18.165 18.515 18.235 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 22.645 17.955 22.715 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 22.365 18.515 22.435 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 25.445 17.955 25.515 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 26.285 18.515 26.355 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 30.485 17.955 30.555 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 29.925 18.515 29.995 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 33.285 17.955 33.355 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 34.125 18.515 34.195 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 38.325 17.955 38.395 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 37.765 18.515 37.835 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 42.245 17.955 42.315 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 41.685 18.515 41.755 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 46.165 17.955 46.235 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 45.885 18.515 45.955 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 50.085 17.955 50.155 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 49.525 18.515 49.595 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 54.005 17.955 54.075 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 53.445 18.515 53.515 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 57.925 17.955 57.995 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 57.645 18.515 57.715 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 61.845 17.955 61.915 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 61.565 18.515 61.635 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 65.765 17.955 65.835 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 65.205 18.515 65.275 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 69.685 17.955 69.755 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 69.405 18.515 69.475 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 73.605 17.955 73.675 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 73.325 18.515 73.395 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 76.405 17.955 76.475 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 77.245 18.515 77.315 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 81.445 17.955 81.515 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 81.165 18.515 81.235 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 84.245 17.955 84.315 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 84.805 18.515 84.875 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 89.285 17.955 89.355 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 88.725 18.515 88.795 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 93.205 17.955 93.275 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 92.925 18.515 92.995 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 97.125 17.955 97.195 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 96.845 18.515 96.915 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 101.045 17.955 101.115 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 100.485 18.515 100.555 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 104.965 17.955 105.035 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 104.685 18.515 104.755 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 108.885 17.955 108.955 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 108.325 18.515 108.395 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 112.805 17.955 112.875 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 112.525 18.515 112.595 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 116.725 17.955 116.795 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 116.445 18.515 116.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 119.525 17.955 119.595 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 120.365 18.515 120.435 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 124.565 17.955 124.635 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 124.285 18.515 124.355 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 147.805 17.955 147.875 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 146.685 18.515 146.755 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 151.725 17.955 151.795 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 150.605 18.515 150.675 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 155.645 17.955 155.715 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 154.525 18.515 154.595 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 159.565 17.955 159.635 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 158.445 18.515 158.515 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 163.485 17.955 163.555 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 162.365 18.515 162.435 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 167.405 17.955 167.475 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 166.285 18.515 166.355 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 171.045 17.955 171.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 170.205 18.515 170.275 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 175.245 17.955 175.315 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 174.125 18.515 174.195 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 178.885 17.955 178.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 179.445 18.515 179.515 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 183.085 17.955 183.155 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 181.965 18.515 182.035 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 186.725 17.955 186.795 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 187.285 18.515 187.355 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 190.925 17.955 190.995 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 189.805 18.515 189.875 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 194.845 17.955 194.915 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 193.725 18.515 193.795 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 198.765 17.955 198.835 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 197.645 18.515 197.715 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 202.685 17.955 202.755 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 201.565 18.515 201.635 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 206.605 17.955 206.675 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 205.485 18.515 205.555 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 210.525 17.955 210.595 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 209.405 18.515 209.475 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 214.445 17.955 214.515 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 213.325 18.515 213.395 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 218.365 17.955 218.435 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 217.245 18.515 217.315 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 222.005 17.955 222.075 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 221.165 18.515 221.235 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 226.205 17.955 226.275 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 225.085 18.515 225.155 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 230.125 17.955 230.195 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 230.405 18.515 230.475 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 234.045 17.955 234.115 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 232.925 18.515 232.995 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 237.965 17.955 238.035 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 236.845 18.515 236.915 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 241.885 17.955 241.955 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 240.765 18.515 240.835 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 245.805 17.955 245.875 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 244.685 18.515 244.755 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 249.725 17.955 249.795 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 248.605 18.515 248.675 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 253.645 17.955 253.715 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 252.525 18.515 252.595 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 257.565 17.955 257.635 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 256.445 18.515 256.515 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 261.485 17.955 261.555 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 260.365 18.515 260.435 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 265.125 17.955 265.195 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 264.285 18.515 264.355 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 269.325 17.955 269.395 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 268.205 18.515 268.275 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p285
    PIN p286
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p287
    PIN p288
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p289
    PIN p290
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p291
    PIN p292
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p293
    PIN p294
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p295
    PIN p296
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 148.085 1.155 148.155 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 152.005 1.155 152.075 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.925 1.155 155.995 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.845 1.155 159.915 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 163.765 1.155 163.835 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 167.685 1.155 167.755 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.605 1.155 171.675 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 175.525 1.155 175.595 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 179.445 1.155 179.515 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 183.365 1.155 183.435 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 187.285 1.155 187.355 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 191.205 1.155 191.275 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 195.125 1.155 195.195 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 199.045 1.155 199.115 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.965 1.155 203.035 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.885 1.155 206.955 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 210.805 1.155 210.875 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 214.725 1.155 214.795 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 218.645 1.155 218.715 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 222.565 1.155 222.635 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 226.485 1.155 226.555 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 230.405 1.155 230.475 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 234.325 1.155 234.395 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 238.245 1.155 238.315 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 242.165 1.155 242.235 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 246.085 1.155 246.155 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 250.005 1.155 250.075 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.925 1.155 253.995 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.845 1.155 257.915 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 261.765 1.155 261.835 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 265.685 1.155 265.755 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 269.605 1.155 269.675 ;
        END
    END p335
    OBS
      LAYER via2 ;
        RECT  0 0 20.16 273.84 ;
      LAYER metal2 ;
        RECT  0 0 20.16 273.84 ;
      LAYER via1 ;
        RECT  0 0 20.16 273.84 ;
      LAYER metal1 ;
        RECT  0 0 20.16 273.84 ;
    END
END fake_macro_newblue1_o330442

MACRO fake_macro_newblue1_o330443
    CLASS BLOCK ;
    SIZE 11.76 BY 268.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.565 9.555 138.635 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.245 1.155 252.315 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.085 1.155 260.155 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.525 1.155 35.595 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.005 1.155 61.075 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.645 1.155 78.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 94.325 1.155 94.395 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.125 1.155 104.195 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.965 1.155 112.035 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.685 1.155 125.755 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.085 1.155 155.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.925 1.155 162.995 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.765 1.155 170.835 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.605 1.155 178.675 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.445 1.155 186.515 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 188.685 1.155 188.755 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.285 1.155 194.355 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 196.525 1.155 196.595 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.125 1.155 202.195 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 204.365 1.155 204.435 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.965 1.155 210.035 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.805 1.155 217.875 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.645 1.155 225.715 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.485 1.155 233.555 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.325 1.155 241.395 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.085 1.155 253.155 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.325 1.155 255.395 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.925 1.155 260.995 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 263.165 1.155 263.235 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 136.605 9.555 136.675 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.325 1.155 136.395 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 131.005 10.115 131.075 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 126.805 10.115 126.875 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.285 9.555 138.355 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.165 1.155 256.235 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.005 1.155 264.075 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 166.285 9.555 166.355 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 120.645 10.115 120.715 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 124.565 10.115 124.635 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 252.245 10.115 252.315 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 256.165 10.115 256.235 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 260.085 10.115 260.155 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 264.005 10.115 264.075 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.805 1.155 252.875 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.645 1.155 260.715 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p265
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER via1 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal1 ;
        RECT  0 0 11.76 268.8 ;
    END
END fake_macro_newblue1_o330443

MACRO fake_macro_newblue1_o330444
    CLASS BLOCK ;
    SIZE 11.76 BY 268.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 124.565 10.115 124.635 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 120.645 10.115 120.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.565 9.555 138.635 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.285 9.555 138.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.525 1.155 35.595 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.005 1.155 61.075 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.645 1.155 78.715 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 94.325 1.155 94.395 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.125 1.155 104.195 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.965 1.155 112.035 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.685 1.155 125.755 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.085 1.155 155.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.925 1.155 162.995 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.765 1.155 170.835 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.605 1.155 178.675 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.445 1.155 186.515 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 188.685 1.155 188.755 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.285 1.155 194.355 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 196.525 1.155 196.595 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.125 1.155 202.195 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 204.365 1.155 204.435 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.965 1.155 210.035 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.805 1.155 217.875 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.645 1.155 225.715 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.485 1.155 233.555 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.325 1.155 241.395 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.085 1.155 253.155 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.325 1.155 255.395 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.925 1.155 260.995 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 263.165 1.155 263.235 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 136.605 9.555 136.675 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.325 1.155 136.395 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 131.005 10.115 131.075 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 126.805 10.115 126.875 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.245 1.155 252.315 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.165 1.155 256.235 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.085 1.155 260.155 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.005 1.155 264.075 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 166.285 9.555 166.355 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 252.245 10.115 252.315 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 256.165 10.115 256.235 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 260.085 10.115 260.155 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 264.005 10.115 264.075 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.805 1.155 252.875 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.645 1.155 260.715 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p265
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER via1 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal1 ;
        RECT  0 0 11.76 268.8 ;
    END
END fake_macro_newblue1_o330444

MACRO fake_macro_newblue1_o330445
    CLASS BLOCK ;
    SIZE 11.76 BY 268.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.565 9.555 138.635 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.285 9.555 138.355 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 166.285 9.555 166.355 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.245 1.155 252.315 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.165 1.155 256.235 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.085 1.155 260.155 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.525 1.155 35.595 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.165 1.155 53.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.005 1.155 61.075 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.645 1.155 78.715 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 94.325 1.155 94.395 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.125 1.155 104.195 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.965 1.155 112.035 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 125.685 1.155 125.755 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 145.565 1.155 145.635 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.085 1.155 155.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.925 1.155 162.995 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.765 1.155 170.835 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.605 1.155 178.675 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.445 1.155 186.515 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 188.685 1.155 188.755 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.285 1.155 194.355 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 196.525 1.155 196.595 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.125 1.155 202.195 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 204.365 1.155 204.435 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.965 1.155 210.035 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.885 1.155 213.955 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.805 1.155 217.875 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.645 1.155 225.715 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.485 1.155 233.555 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.325 1.155 241.395 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.245 1.155 245.315 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.485 1.155 247.555 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.085 1.155 253.155 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.325 1.155 255.395 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.925 1.155 260.995 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 263.165 1.155 263.235 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 131.005 10.115 131.075 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 126.805 10.115 126.875 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 136.605 9.555 136.675 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.325 1.155 136.395 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.005 1.155 264.075 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 18.725 10.115 18.795 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 22.645 10.115 22.715 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 26.565 10.115 26.635 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 30.485 10.115 30.555 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 34.405 10.115 34.475 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 38.325 10.115 38.395 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 42.245 10.115 42.315 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 46.165 10.115 46.235 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 50.085 10.115 50.155 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 54.005 10.115 54.075 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 57.925 10.115 57.995 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 61.845 10.115 61.915 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 65.765 10.115 65.835 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 69.685 10.115 69.755 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 73.605 10.115 73.675 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 77.525 10.115 77.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 81.445 10.115 81.515 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 85.365 10.115 85.435 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 89.285 10.115 89.355 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 93.205 10.115 93.275 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 97.125 10.115 97.195 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 101.045 10.115 101.115 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 104.965 10.115 105.035 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 108.885 10.115 108.955 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 112.805 10.115 112.875 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 116.725 10.115 116.795 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 120.645 10.115 120.715 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 124.565 10.115 124.635 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 142.485 10.115 142.555 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 146.405 10.115 146.475 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 150.325 10.115 150.395 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 158.165 10.115 158.235 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 162.085 10.115 162.155 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 166.005 10.115 166.075 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 169.925 10.115 169.995 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 173.845 10.115 173.915 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 177.765 10.115 177.835 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 181.685 10.115 181.755 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 185.605 10.115 185.675 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 189.525 10.115 189.595 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 193.445 10.115 193.515 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 197.365 10.115 197.435 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 201.285 10.115 201.355 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 205.205 10.115 205.275 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 209.125 10.115 209.195 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 213.045 10.115 213.115 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 216.965 10.115 217.035 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 220.885 10.115 220.955 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 224.805 10.115 224.875 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 228.725 10.115 228.795 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 232.645 10.115 232.715 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 236.565 10.115 236.635 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 240.485 10.115 240.555 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 244.405 10.115 244.475 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 248.325 10.115 248.395 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 252.245 10.115 252.315 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 256.165 10.115 256.235 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 260.085 10.115 260.155 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 264.005 10.115 264.075 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.805 1.155 252.875 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.645 1.155 260.715 ;
        END
    END p265
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal2 ;
        RECT  0 0 11.76 268.8 ;
      LAYER via1 ;
        RECT  0 0 11.76 268.8 ;
      LAYER metal1 ;
        RECT  0 0 11.76 268.8 ;
    END
END fake_macro_newblue1_o330445

MACRO fake_macro_newblue1_o330446
    CLASS BLOCK ;
    SIZE 15.68 BY 142.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.885 13.475 73.955 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 83.685 14.035 83.755 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 79.765 14.035 79.835 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.805 1.155 21.875 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.645 1.155 127.715 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.285 1.155 110.355 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 68.285 14.035 68.355 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 64.085 14.035 64.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 71.365 1.155 71.435 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.245 1.155 70.315 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.845 13.475 75.915 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.565 13.475 75.635 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.845 1.155 82.915 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.765 1.155 79.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.685 1.155 83.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 103.565 13.475 103.635 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.325 1.155 80.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.245 1.155 84.315 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p139
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER via1 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal1 ;
        RECT  0 0 15.68 142.8 ;
    END
END fake_macro_newblue1_o330446

MACRO fake_macro_newblue1_o330447
    CLASS BLOCK ;
    SIZE 15.68 BY 142.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.885 13.475 73.955 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 107.205 14.035 107.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 103.285 14.035 103.355 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 99.365 14.035 99.435 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 95.445 14.035 95.515 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 91.525 14.035 91.595 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 87.605 14.035 87.675 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 83.685 14.035 83.755 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 79.765 14.035 79.835 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 61.845 14.035 61.915 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 138.565 14.035 138.635 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 134.645 14.035 134.715 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 130.725 14.035 130.795 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 126.805 14.035 126.875 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 122.885 14.035 122.955 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 118.965 14.035 119.035 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 115.045 14.035 115.115 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 111.125 14.035 111.195 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 71.365 1.155 71.435 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 38.325 14.035 38.395 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 34.405 14.035 34.475 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 30.485 14.035 30.555 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 54.005 14.035 54.075 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 22.645 14.035 22.715 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 18.725 14.035 18.795 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 57.925 14.035 57.995 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 50.085 14.035 50.155 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 46.165 14.035 46.235 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 42.245 14.035 42.315 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 26.565 14.035 26.635 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.845 13.475 75.915 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 75.565 13.475 75.635 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 103.565 13.475 103.635 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.845 1.155 82.915 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.645 1.155 127.715 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.285 1.155 110.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.685 1.155 76.755 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 68.285 14.035 68.355 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 64.085 14.035 64.155 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.245 1.155 70.315 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.805 1.155 21.875 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.765 1.155 79.835 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.685 1.155 83.755 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.325 1.155 80.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.245 1.155 84.315 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.165 1.155 88.235 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.085 1.155 92.155 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.005 1.155 96.075 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.925 1.155 99.995 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.845 1.155 103.915 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.765 1.155 107.835 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.685 1.155 111.755 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.605 1.155 115.675 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.525 1.155 119.595 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.445 1.155 123.515 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.365 1.155 127.435 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.285 1.155 131.355 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.205 1.155 135.275 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.125 1.155 139.195 ;
        END
    END p139
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal2 ;
        RECT  0 0 15.68 142.8 ;
      LAYER via1 ;
        RECT  0 0 15.68 142.8 ;
      LAYER metal1 ;
        RECT  0 0 15.68 142.8 ;
    END
END fake_macro_newblue1_o330447

MACRO fake_macro_newblue1_o330448
    CLASS BLOCK ;
    SIZE 11.76 BY 48.72 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.645 1.155 43.715 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.725 1.155 39.795 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.885 1.155 31.955 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 13.965 1.155 14.035 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.125 1.155 6.195 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 28.805 9.555 28.875 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 28.525 9.555 28.595 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 48.405 9.555 48.475 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 26.845 9.555 26.915 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 21.245 10.115 21.315 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 17.045 10.115 17.115 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 32.725 1.155 32.795 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 36.645 1.155 36.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 40.565 1.155 40.635 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 44.485 1.155 44.555 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 32.725 10.115 32.795 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 36.645 10.115 36.715 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 40.565 10.115 40.635 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 44.485 10.115 44.555 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.285 1.155 33.355 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.205 1.155 37.275 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.125 1.155 41.195 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.045 1.155 45.115 ;
        END
    END p41
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 48.72 ;
      LAYER metal2 ;
        RECT  0 0 11.76 48.72 ;
      LAYER via1 ;
        RECT  0 0 11.76 48.72 ;
      LAYER metal1 ;
        RECT  0 0 11.76 48.72 ;
    END
END fake_macro_newblue1_o330448

MACRO fake_macro_newblue1_o330449
    CLASS BLOCK ;
    SIZE 15.68 BY 48.72 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 28.805 13.475 28.875 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 24.325 1.155 24.395 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.845 13.475 26.915 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 21.245 14.035 21.315 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 17.045 14.035 17.115 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.205 1.155 23.275 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 28.525 13.475 28.595 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 32.725 1.155 32.795 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 36.645 1.155 36.715 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 40.565 1.155 40.635 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 44.485 1.155 44.555 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 48.405 13.475 48.475 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 32.725 14.035 32.795 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 36.645 14.035 36.715 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 40.565 14.035 40.635 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 44.485 14.035 44.555 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.285 1.155 33.355 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.205 1.155 37.275 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.125 1.155 41.195 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.045 1.155 45.115 ;
        END
    END p43
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 48.72 ;
      LAYER metal2 ;
        RECT  0 0 15.68 48.72 ;
      LAYER via1 ;
        RECT  0 0 15.68 48.72 ;
      LAYER metal1 ;
        RECT  0 0 15.68 48.72 ;
    END
END fake_macro_newblue1_o330449

MACRO fake_macro_newblue1_o330450
    CLASS BLOCK ;
    SIZE 15.68 BY 48.72 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.845 13.475 26.915 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 28.805 13.475 28.875 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 21.245 14.035 21.315 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 17.045 14.035 17.115 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 24.325 1.155 24.395 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.205 1.155 23.275 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 48.405 13.475 48.475 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 28.525 13.475 28.595 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 32.725 1.155 32.795 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 36.645 1.155 36.715 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 40.565 1.155 40.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 44.485 1.155 44.555 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 32.725 14.035 32.795 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 36.645 14.035 36.715 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 40.565 14.035 40.635 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 44.485 14.035 44.555 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.285 1.155 33.355 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.205 1.155 37.275 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.125 1.155 41.195 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.045 1.155 45.115 ;
        END
    END p43
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 48.72 ;
      LAYER metal2 ;
        RECT  0 0 15.68 48.72 ;
      LAYER via1 ;
        RECT  0 0 15.68 48.72 ;
      LAYER metal1 ;
        RECT  0 0 15.68 48.72 ;
    END
END fake_macro_newblue1_o330450

MACRO fake_macro_newblue1_o330451
    CLASS BLOCK ;
    SIZE 11.76 BY 48.72 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.045 1.155 45.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.645 1.155 43.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.725 1.155 39.795 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.885 1.155 31.955 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 13.965 1.155 14.035 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.045 1.155 10.115 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.125 1.155 6.195 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.205 1.155 2.275 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 28.805 9.555 28.875 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 48.405 9.555 48.475 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 26.845 9.555 26.915 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 21.245 10.115 21.315 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 17.045 10.115 17.115 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 28.525 9.555 28.595 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 32.725 1.155 32.795 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 36.645 1.155 36.715 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 40.565 1.155 40.635 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 44.485 1.155 44.555 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 3.045 10.115 3.115 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 6.965 10.115 7.035 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 10.885 10.115 10.955 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 14.805 10.115 14.875 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 32.725 10.115 32.795 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 36.645 10.115 36.715 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 40.565 10.115 40.635 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 44.485 10.115 44.555 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.285 1.155 33.355 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.205 1.155 37.275 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.125 1.155 41.195 ;
        END
    END p41
    OBS
      LAYER via2 ;
        RECT  0 0 11.76 48.72 ;
      LAYER metal2 ;
        RECT  0 0 11.76 48.72 ;
      LAYER via1 ;
        RECT  0 0 11.76 48.72 ;
      LAYER metal1 ;
        RECT  0 0 11.76 48.72 ;
    END
END fake_macro_newblue1_o330451

MACRO fake_macro_newblue1_o330452
    CLASS BLOCK ;
    SIZE 15.68 BY 48.72 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 24.325 1.155 24.395 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.845 13.475 26.915 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 28.805 13.475 28.875 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 21.245 14.035 21.315 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 17.045 14.035 17.115 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.205 1.155 23.275 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 28.525 13.475 28.595 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 32.725 1.155 32.795 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 36.645 1.155 36.715 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 40.565 1.155 40.635 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 44.485 1.155 44.555 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 48.405 13.475 48.475 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 32.725 14.035 32.795 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 36.645 14.035 36.715 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 40.565 14.035 40.635 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 44.485 14.035 44.555 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.285 1.155 33.355 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.205 1.155 37.275 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.125 1.155 41.195 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.045 1.155 45.115 ;
        END
    END p43
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 48.72 ;
      LAYER metal2 ;
        RECT  0 0 15.68 48.72 ;
      LAYER via1 ;
        RECT  0 0 15.68 48.72 ;
      LAYER metal1 ;
        RECT  0 0 15.68 48.72 ;
    END
END fake_macro_newblue1_o330452

MACRO fake_macro_newblue1_o330453
    CLASS BLOCK ;
    SIZE 15.68 BY 48.72 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.325 1.155 45.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.485 1.155 37.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.845 13.475 26.915 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 28.805 13.475 28.875 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 28.525 13.475 28.595 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.645 1.155 29.715 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 21.245 14.035 21.315 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 17.045 14.035 17.115 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 24.325 1.155 24.395 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.205 1.155 23.275 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 32.725 1.155 32.795 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 36.645 1.155 36.715 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 40.565 1.155 40.635 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 44.485 1.155 44.555 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 48.405 13.475 48.475 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 3.045 14.035 3.115 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 6.965 14.035 7.035 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 10.885 14.035 10.955 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 14.805 14.035 14.875 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 32.725 14.035 32.795 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 36.645 14.035 36.715 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 40.565 14.035 40.635 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 44.485 14.035 44.555 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.285 1.155 33.355 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.205 1.155 37.275 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.125 1.155 41.195 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.045 1.155 45.115 ;
        END
    END p43
    OBS
      LAYER via2 ;
        RECT  0 0 15.68 48.72 ;
      LAYER metal2 ;
        RECT  0 0 15.68 48.72 ;
      LAYER via1 ;
        RECT  0 0 15.68 48.72 ;
      LAYER metal1 ;
        RECT  0 0 15.68 48.72 ;
    END
END fake_macro_newblue1_o330453

MACRO fake_macro_newblue1_o330454
    CLASS BLOCK ;
    SIZE 23.52 BY 268.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 138.565 21.315 138.635 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.245 1.155 252.315 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.165 1.155 256.235 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.085 1.155 260.155 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.005 1.155 264.075 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.125 1.155 6.195 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.405 1.155 41.475 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.085 1.155 57.155 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.645 1.155 78.715 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 98.245 1.155 98.315 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.845 1.155 117.915 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.765 1.155 121.835 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 141.645 1.155 141.715 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.245 1.155 147.315 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.165 1.155 151.235 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.925 1.155 162.995 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.765 1.155 170.835 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.605 1.155 178.675 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.605 1.155 192.675 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.125 1.155 202.195 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.285 1.155 208.355 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 212.205 1.155 212.275 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.805 1.155 217.875 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.645 1.155 225.715 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.485 1.155 233.555 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.325 1.155 241.395 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 243.565 1.155 243.635 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 249.165 1.155 249.235 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.085 1.155 253.155 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.005 1.155 257.075 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 259.245 1.155 259.315 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.845 1.155 264.915 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.605 21.315 136.675 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.045 1.155 136.115 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 131.005 21.875 131.075 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 126.805 21.875 126.875 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.085 1.155 134.155 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.965 1.155 133.035 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.085 2.275 134.155 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 132.965 2.275 133.035 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 138.285 21.315 138.355 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 166.285 21.315 166.355 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 3.045 21.875 3.115 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 6.965 21.875 7.035 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 10.885 21.875 10.955 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 14.805 21.875 14.875 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 18.725 21.875 18.795 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 22.645 21.875 22.715 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 26.565 21.875 26.635 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 30.485 21.875 30.555 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 34.405 21.875 34.475 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 38.325 21.875 38.395 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 42.245 21.875 42.315 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 46.165 21.875 46.235 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 50.085 21.875 50.155 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 54.005 21.875 54.075 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 57.925 21.875 57.995 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 61.845 21.875 61.915 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 65.765 21.875 65.835 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 69.685 21.875 69.755 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 73.605 21.875 73.675 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 77.525 21.875 77.595 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 81.445 21.875 81.515 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 85.365 21.875 85.435 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 89.285 21.875 89.355 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 93.205 21.875 93.275 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 97.125 21.875 97.195 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 101.045 21.875 101.115 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 104.965 21.875 105.035 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 108.885 21.875 108.955 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 112.805 21.875 112.875 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 116.725 21.875 116.795 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 120.645 21.875 120.715 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 124.565 21.875 124.635 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 142.485 21.875 142.555 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 146.405 21.875 146.475 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 150.325 21.875 150.395 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 154.245 21.875 154.315 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 158.165 21.875 158.235 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 162.085 21.875 162.155 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 166.005 21.875 166.075 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 169.925 21.875 169.995 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 173.845 21.875 173.915 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 177.765 21.875 177.835 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 181.685 21.875 181.755 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 185.605 21.875 185.675 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 189.525 21.875 189.595 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 193.445 21.875 193.515 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 197.365 21.875 197.435 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 201.285 21.875 201.355 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 205.205 21.875 205.275 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 209.125 21.875 209.195 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 213.045 21.875 213.115 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 216.965 21.875 217.035 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 220.885 21.875 220.955 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 224.805 21.875 224.875 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 228.725 21.875 228.795 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 232.645 21.875 232.715 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 236.565 21.875 236.635 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 240.485 21.875 240.555 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 244.405 21.875 244.475 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 248.325 21.875 248.395 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 252.245 21.875 252.315 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 256.165 21.875 256.235 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 260.085 21.875 260.155 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 264.005 21.875 264.075 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.805 1.155 252.875 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.645 1.155 260.715 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p269
    OBS
      LAYER via2 ;
        RECT  0 0 23.52 268.8 ;
      LAYER metal2 ;
        RECT  0 0 23.52 268.8 ;
      LAYER via1 ;
        RECT  0 0 23.52 268.8 ;
      LAYER metal1 ;
        RECT  0 0 23.52 268.8 ;
    END
END fake_macro_newblue1_o330454

MACRO fake_macro_newblue1_o330455
    CLASS BLOCK ;
    SIZE 71.96 BY 307.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 303.765 1.155 303.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 297.885 2.275 297.955 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 290.045 2.275 290.115 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 282.205 2.275 282.275 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.365 2.275 274.435 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.525 2.275 266.595 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.685 2.275 258.755 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.845 2.275 250.915 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 243.005 2.275 243.075 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 235.165 2.275 235.235 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.325 2.275 227.395 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.485 2.275 219.555 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.645 2.275 211.715 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.805 2.275 203.875 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.965 2.275 196.035 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 188.125 2.275 188.195 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.285 2.275 180.355 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.445 2.275 172.515 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.605 2.275 164.675 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.765 2.275 156.835 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 135.205 2.275 135.275 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.365 2.275 127.435 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.525 2.275 119.595 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.685 2.275 111.755 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.845 2.275 103.915 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 96.005 2.275 96.075 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 88.165 2.275 88.235 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.325 2.275 80.395 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.485 2.275 72.555 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.645 2.275 64.715 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.805 2.275 56.875 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.965 2.275 49.035 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 41.125 2.275 41.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.285 2.275 33.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.445 2.275 25.515 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.605 2.275 17.675 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.765 2.275 9.835 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.925 2.275 1.995 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 149.765 3.955 149.835 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.765 2.275 149.835 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 149.765 1.155 149.835 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.445 1.155 151.515 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 152.005 1.155 152.075 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.365 69.475 148.435 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.285 69.475 152.355 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 144.445 1.155 144.515 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 170.205 69.475 170.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.245 1.155 147.315 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.645 3.955 148.715 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 154.245 69.475 154.315 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 154.525 70.035 154.595 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.885 1.155 3.955 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.165 1.155 11.235 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.005 1.155 19.075 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.845 1.155 26.915 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.245 1.155 35.315 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.525 1.155 42.595 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.925 1.155 50.995 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.765 1.155 58.835 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.045 1.155 66.115 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.445 1.155 74.515 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.725 1.155 81.795 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.125 1.155 90.195 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.405 1.155 97.475 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.245 1.155 105.315 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.085 1.155 113.155 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.485 1.155 121.555 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.765 1.155 128.835 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.165 1.155 137.235 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 302.085 1.155 302.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.405 69.475 153.475 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.085 1.155 155.155 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 6.965 70.595 7.035 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 14.805 70.595 14.875 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 23.765 70.595 23.835 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 30.485 70.595 30.555 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 38.325 70.595 38.395 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 46.165 70.595 46.235 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 54.005 70.595 54.075 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 62.965 70.595 63.035 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 69.685 70.595 69.755 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 77.525 70.595 77.595 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 86.485 70.595 86.555 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 93.205 70.595 93.275 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 101.045 70.595 101.115 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 108.885 70.595 108.955 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 116.725 70.595 116.795 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 125.685 70.595 125.755 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 132.405 70.595 132.475 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 140.245 70.595 140.315 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 157.045 70.595 157.115 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 164.885 70.595 164.955 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 173.845 70.595 173.915 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 180.565 70.595 180.635 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 189.525 70.595 189.595 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 197.365 70.595 197.435 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 205.205 70.595 205.275 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 211.925 70.595 211.995 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 219.765 70.595 219.835 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 227.605 70.595 227.675 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 235.445 70.595 235.515 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 243.285 70.595 243.355 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 251.125 70.595 251.195 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 260.085 70.595 260.155 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 266.805 70.595 266.875 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 274.645 70.595 274.715 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 283.605 70.595 283.675 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 290.325 70.595 290.395 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 298.165 70.595 298.235 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 272.405 1.155 272.475 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 280.245 1.155 280.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 288.085 1.155 288.155 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 295.925 1.155 295.995 ;
        END
    END p167
    OBS
      LAYER via2 ;
        RECT  0 0 72.1 307.44 ;
      LAYER metal2 ;
        RECT  0 0 72.1 307.44 ;
      LAYER via1 ;
        RECT  0 0 72.1 307.44 ;
      LAYER metal1 ;
        RECT  0 0 72.1 307.44 ;
    END
END fake_macro_newblue1_o330455

MACRO fake_macro_newblue1_o330456
    CLASS BLOCK ;
    SIZE 70.56 BY 146.16 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 51.205 1.155 51.275 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.845 1.155 82.915 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.445 1.155 102.515 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.365 1.155 106.435 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.285 1.155 110.355 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.885 1.155 129.955 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 133.805 1.155 133.875 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.725 1.155 137.795 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.605 1.155 143.675 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.765 1.155 142.835 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.925 1.155 134.995 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.005 1.155 131.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.245 1.155 119.315 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.805 1.155 91.875 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.885 1.155 87.955 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.685 1.155 34.755 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.925 1.155 22.995 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.165 1.155 11.235 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.605 1.155 80.675 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.365 1.155 50.435 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.965 68.355 70.035 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 71.925 68.355 71.995 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.205 1.155 72.275 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 77.525 68.915 77.595 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 72.765 1.155 72.835 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 81.725 68.915 81.795 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.445 1.155 74.515 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 75.565 1.155 75.635 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 73.325 1.715 73.395 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 75.565 1.715 75.635 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 74.445 3.395 74.515 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 75.565 3.395 75.635 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 74.445 1.715 74.515 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 76.685 1.715 76.755 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 97.685 68.355 97.755 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 70.245 68.355 70.315 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.845 1.155 138.915 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.085 1.155 127.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.165 1.155 123.235 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.325 1.155 115.395 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.405 1.155 111.475 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.485 1.155 107.555 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.565 1.155 103.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.645 1.155 99.715 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.725 1.155 95.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.965 1.155 84.035 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.045 1.155 66.115 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.125 1.155 62.195 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.285 1.155 54.355 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.445 1.155 46.515 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.525 1.155 42.595 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.605 1.155 38.675 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.765 1.155 30.835 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.845 1.155 26.915 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.005 1.155 19.075 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.085 1.155 15.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.245 1.155 7.315 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.325 1.155 3.395 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.765 68.915 142.835 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 138.845 68.915 138.915 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 134.925 68.915 134.995 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 131.005 68.915 131.075 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 127.085 68.915 127.155 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 123.165 68.915 123.235 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 119.245 68.915 119.315 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 115.325 68.915 115.395 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 111.405 68.915 111.475 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 107.485 68.915 107.555 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 103.565 68.915 103.635 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 99.645 68.915 99.715 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 95.725 68.915 95.795 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 91.805 68.915 91.875 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 87.885 68.915 87.955 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 83.965 68.915 84.035 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 66.045 68.915 66.115 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 62.125 68.915 62.195 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 58.205 68.915 58.275 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 54.285 68.915 54.355 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 50.365 68.915 50.435 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 46.445 68.915 46.515 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 42.525 68.915 42.595 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 38.605 68.915 38.675 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 34.685 68.915 34.755 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 30.765 68.915 30.835 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 26.845 68.915 26.915 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 22.925 68.915 22.995 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 19.005 68.915 19.075 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 15.085 68.915 15.155 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 11.165 68.915 11.235 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 7.245 68.915 7.315 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 3.325 68.915 3.395 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.485 1.155 135.555 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 131.565 1.155 131.635 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.645 1.155 127.715 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 119.805 1.155 119.875 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.965 1.155 112.035 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.045 1.155 108.115 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.125 1.155 104.195 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.205 1.155 100.275 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.285 1.155 96.355 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.445 1.155 88.515 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.525 1.155 84.595 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.485 1.155 65.555 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.565 1.155 61.635 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.645 1.155 57.715 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.725 1.155 53.795 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.805 1.155 49.875 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.885 1.155 45.955 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.965 1.155 42.035 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.045 1.155 38.115 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.125 1.155 34.195 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.205 1.155 30.275 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.285 1.155 26.355 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.365 1.155 22.435 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.445 1.155 18.515 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.525 1.155 14.595 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.605 1.155 10.675 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.685 1.155 6.755 ;
        END
    END p149
    OBS
      LAYER via2 ;
        RECT  0 0 70.56 146.16 ;
      LAYER metal2 ;
        RECT  0 0 70.56 146.16 ;
      LAYER via1 ;
        RECT  0 0 70.56 146.16 ;
      LAYER metal1 ;
        RECT  0 0 70.56 146.16 ;
    END
END fake_macro_newblue1_o330456

MACRO fake_macro_newblue1_o330457
    CLASS BLOCK ;
    SIZE 71.96 BY 307.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 303.765 1.155 303.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 297.885 2.275 297.955 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 290.045 2.275 290.115 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 282.205 2.275 282.275 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.365 2.275 274.435 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.525 2.275 266.595 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.685 2.275 258.755 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.845 2.275 250.915 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 243.005 2.275 243.075 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 235.165 2.275 235.235 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.325 2.275 227.395 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.485 2.275 219.555 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.645 2.275 211.715 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.805 2.275 203.875 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.965 2.275 196.035 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 188.125 2.275 188.195 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.285 2.275 180.355 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.445 2.275 172.515 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.605 2.275 164.675 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.765 2.275 156.835 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 135.205 2.275 135.275 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.365 2.275 127.435 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.525 2.275 119.595 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.685 2.275 111.755 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.845 2.275 103.915 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 96.005 2.275 96.075 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 88.165 2.275 88.235 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.325 2.275 80.395 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.485 2.275 72.555 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.645 2.275 64.715 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.805 2.275 56.875 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.965 2.275 49.035 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 41.125 2.275 41.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.285 2.275 33.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.445 2.275 25.515 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.605 2.275 17.675 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.765 2.275 9.835 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.925 2.275 1.995 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.405 69.475 153.475 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.845 1.155 26.915 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.645 3.955 148.715 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 144.445 1.155 144.515 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 154.245 69.475 154.315 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 181.965 69.475 182.035 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.525 1.155 42.595 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.725 1.155 81.795 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.125 1.155 90.195 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.405 1.155 97.475 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.485 1.155 121.555 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 137.165 1.155 137.235 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 302.085 1.155 302.155 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.245 1.155 35.315 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 298.165 70.595 298.235 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 260.085 70.595 260.155 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 251.125 70.595 251.195 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 243.285 70.595 243.355 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 235.445 70.595 235.515 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 227.605 70.595 227.675 ;
        END
    END p68
    PIN p69
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 219.765 70.595 219.835 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 211.925 70.595 211.995 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 205.205 70.595 205.275 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 197.365 70.595 197.435 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 189.525 70.595 189.595 ;
        END
    END p73
    PIN p74
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 180.565 70.595 180.635 ;
        END
    END p74
    PIN p75
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 173.845 70.595 173.915 ;
        END
    END p75
    PIN p76
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 164.885 70.595 164.955 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 157.045 70.595 157.115 ;
        END
    END p77
    PIN p78
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 140.245 70.595 140.315 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 132.405 70.595 132.475 ;
        END
    END p79
    PIN p80
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 125.685 70.595 125.755 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 116.725 70.595 116.795 ;
        END
    END p81
    PIN p82
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 108.885 70.595 108.955 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 101.045 70.595 101.115 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 93.205 70.595 93.275 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 86.485 70.595 86.555 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 77.525 70.595 77.595 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 69.685 70.595 69.755 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 62.965 70.595 63.035 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 54.005 70.595 54.075 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 46.165 70.595 46.235 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 38.325 70.595 38.395 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 30.485 70.595 30.555 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 23.765 70.595 23.835 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 14.805 70.595 14.875 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 6.965 70.595 7.035 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 290.325 70.595 290.395 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 283.605 70.595 283.675 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 274.645 70.595 274.715 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 266.805 70.595 266.875 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.285 69.475 152.355 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.365 69.475 148.435 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 152.005 1.155 152.075 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.445 1.155 151.515 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.965 69.475 154.035 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 149.765 1.155 149.835 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.245 1.155 147.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.765 2.275 149.835 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 149.765 3.955 149.835 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.885 1.155 3.955 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.165 1.155 11.235 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.005 1.155 19.075 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.925 1.155 50.995 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.765 1.155 58.835 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.045 1.155 66.115 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.445 1.155 74.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.245 1.155 105.315 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.085 1.155 113.155 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 128.765 1.155 128.835 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.445 1.155 200.515 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.805 1.155 231.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.085 1.155 155.155 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 272.405 1.155 272.475 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 280.245 1.155 280.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 288.085 1.155 288.155 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 295.925 1.155 295.995 ;
        END
    END p167
    OBS
      LAYER via2 ;
        RECT  0 0 72.1 307.44 ;
      LAYER metal2 ;
        RECT  0 0 72.1 307.44 ;
      LAYER via1 ;
        RECT  0 0 72.1 307.44 ;
      LAYER metal1 ;
        RECT  0 0 72.1 307.44 ;
    END
END fake_macro_newblue1_o330457

MACRO fake_macro_newblue1_o330458
    CLASS BLOCK ;
    SIZE 70.56 BY 146.16 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 143.045 68.915 143.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 141.645 68.915 141.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 139.405 68.915 139.475 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 135.485 68.915 135.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 131.565 68.915 131.635 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 125.965 68.915 126.035 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 122.045 68.915 122.115 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 118.125 68.915 118.195 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 114.205 68.915 114.275 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 111.965 68.915 112.035 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 108.045 68.915 108.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 104.125 68.915 104.195 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 98.525 68.915 98.595 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 94.605 68.915 94.675 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 90.685 68.915 90.755 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 86.765 68.915 86.835 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 84.525 68.915 84.595 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 80.605 68.915 80.675 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 62.965 68.915 63.035 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 57.085 68.915 57.155 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 53.165 68.915 53.235 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 49.245 68.915 49.315 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 45.325 68.915 45.395 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 43.365 68.915 43.435 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 39.445 68.915 39.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 35.525 68.915 35.595 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 29.645 68.915 29.715 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 25.725 68.915 25.795 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 21.805 68.915 21.875 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 17.885 68.915 17.955 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 15.925 68.915 15.995 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 12.005 68.915 12.075 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 8.085 68.915 8.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 2.205 68.915 2.275 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 71.365 68.355 71.435 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 71.365 66.675 71.435 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 72.485 68.355 72.555 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 71.365 68.915 71.435 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 73.045 68.915 73.115 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 73.605 68.915 73.675 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 3.045 68.915 3.115 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 6.965 68.915 7.035 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 10.885 68.915 10.955 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 18.725 68.915 18.795 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 22.645 68.915 22.715 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 26.565 68.915 26.635 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 30.485 68.915 30.555 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 34.405 68.915 34.475 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 38.325 68.915 38.395 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 42.245 68.915 42.315 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 46.165 68.915 46.235 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 50.085 68.915 50.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 54.005 68.915 54.075 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 57.925 68.915 57.995 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 61.845 68.915 61.915 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 83.685 68.915 83.755 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 87.605 68.915 87.675 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 91.525 68.915 91.595 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 95.445 68.915 95.515 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 99.365 68.915 99.435 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 103.285 68.915 103.355 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 107.205 68.915 107.275 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 111.125 68.915 111.195 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 115.045 68.915 115.115 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 118.965 68.915 119.035 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 122.885 68.915 122.955 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 126.805 68.915 126.875 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 134.645 68.915 134.715 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 75.845 1.715 75.915 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 75.565 1.715 75.635 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 73.885 1.715 73.955 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 65.205 68.915 65.275 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 68.285 1.155 68.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.085 1.155 64.155 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 70.245 68.915 70.315 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 70.245 68.355 70.315 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 70.245 66.675 70.315 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.125 68.355 69.195 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 103.565 1.715 103.635 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 14.805 68.915 14.875 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 79.765 68.915 79.835 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 130.725 68.915 130.795 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 138.565 68.915 138.635 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.485 68.915 142.555 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 76.685 68.915 76.755 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 79.765 1.155 79.835 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 83.685 1.155 83.755 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 87.605 1.155 87.675 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 91.525 1.155 91.595 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 95.445 1.155 95.515 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 99.365 1.155 99.435 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 103.285 1.155 103.355 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 107.205 1.155 107.275 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 111.125 1.155 111.195 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.045 1.155 115.115 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 118.965 1.155 119.035 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 122.885 1.155 122.955 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 126.805 1.155 126.875 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 130.725 1.155 130.795 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.645 1.155 134.715 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 2.485 68.915 2.555 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 6.405 68.915 6.475 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 10.325 68.915 10.395 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 14.245 68.915 14.315 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 18.165 68.915 18.235 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 22.085 68.915 22.155 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 26.005 68.915 26.075 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 29.925 68.915 29.995 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 33.845 68.915 33.915 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 37.765 68.915 37.835 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 41.685 68.915 41.755 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 45.605 68.915 45.675 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 49.525 68.915 49.595 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 53.445 68.915 53.515 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 57.365 68.915 57.435 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 61.285 68.915 61.355 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 80.325 68.915 80.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 84.245 68.915 84.315 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 88.165 68.915 88.235 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 92.085 68.915 92.155 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 96.005 68.915 96.075 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 99.925 68.915 99.995 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 103.845 68.915 103.915 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 107.765 68.915 107.835 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 111.685 68.915 111.755 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 115.605 68.915 115.675 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 119.525 68.915 119.595 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 123.445 68.915 123.515 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 127.365 68.915 127.435 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 131.285 68.915 131.355 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 135.205 68.915 135.275 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 139.125 68.915 139.195 ;
        END
    END p149
    OBS
      LAYER via2 ;
        RECT  0 0 70.56 146.16 ;
      LAYER metal2 ;
        RECT  0 0 70.56 146.16 ;
      LAYER via1 ;
        RECT  0 0 70.56 146.16 ;
      LAYER metal1 ;
        RECT  0 0 70.56 146.16 ;
    END
END fake_macro_newblue1_o330458

MACRO fake_macro_newblue1_o330459
    CLASS BLOCK ;
    SIZE 39.2 BY 268.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.645 1.155 260.715 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.565 1.155 264.635 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 138.565 36.995 138.635 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 142.485 1.155 142.555 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.405 1.155 146.475 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.325 1.155 150.395 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.245 1.155 154.315 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.165 1.155 158.235 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.085 1.155 162.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.005 1.155 166.075 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 169.925 1.155 169.995 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 173.845 1.155 173.915 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 177.765 1.155 177.835 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 181.685 1.155 181.755 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 185.605 1.155 185.675 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 189.525 1.155 189.595 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 193.445 1.155 193.515 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.365 1.155 197.435 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.285 1.155 201.355 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.205 1.155 205.275 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.125 1.155 209.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.045 1.155 213.115 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 216.965 1.155 217.035 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 220.885 1.155 220.955 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 224.805 1.155 224.875 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 228.725 1.155 228.795 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 232.645 1.155 232.715 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 236.565 1.155 236.635 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 240.485 1.155 240.555 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.405 1.155 244.475 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.325 1.155 248.395 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.245 1.155 252.315 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.165 1.155 256.235 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.085 1.155 260.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.005 1.155 264.075 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 4.165 1.155 4.235 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.125 1.155 6.195 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 12.005 1.155 12.075 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 15.925 1.155 15.995 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.845 1.155 19.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.685 1.155 27.755 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 31.605 1.155 31.675 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.565 1.155 33.635 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 39.445 1.155 39.515 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 47.285 1.155 47.355 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.245 1.155 49.315 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 55.125 1.155 55.195 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 59.045 1.155 59.115 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 62.965 1.155 63.035 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 64.925 1.155 64.995 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 70.805 1.155 70.875 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.725 1.155 74.795 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.645 1.155 78.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.565 1.155 82.635 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 86.485 1.155 86.555 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 90.405 1.155 90.475 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.365 1.155 92.435 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 98.245 1.155 98.315 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 102.165 1.155 102.235 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 106.085 1.155 106.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 110.005 1.155 110.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.925 1.155 113.995 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 115.885 1.155 115.955 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.765 1.155 121.835 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 123.725 1.155 123.795 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.325 1.155 143.395 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.245 1.155 147.315 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 149.485 1.155 149.555 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 153.405 1.155 153.475 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.005 1.155 159.075 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.925 1.155 162.995 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.845 1.155 166.915 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.765 1.155 170.835 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.685 1.155 174.755 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.605 1.155 178.675 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.525 1.155 182.595 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.765 1.155 184.835 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.365 1.155 190.435 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.285 1.155 194.355 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.205 1.155 198.275 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.125 1.155 202.195 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.045 1.155 206.115 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.965 1.155 210.035 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 212.205 1.155 212.275 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.805 1.155 217.875 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.725 1.155 221.795 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.645 1.155 225.715 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.565 1.155 229.635 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.485 1.155 233.555 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.405 1.155 237.475 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.325 1.155 241.395 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 243.565 1.155 243.635 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 249.165 1.155 249.235 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 251.405 1.155 251.475 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.005 1.155 257.075 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 260.925 1.155 260.995 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 264.845 1.155 264.915 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 139.405 1.155 139.475 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 138.285 36.995 138.355 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 166.285 36.995 166.355 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 136.605 36.995 136.675 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.925 1.155 127.995 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.325 1.155 136.395 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 131.005 37.555 131.075 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 135.765 1.155 135.835 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 126.805 37.555 126.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 134.085 1.155 134.155 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.965 1.155 133.035 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 134.085 1.715 134.155 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 132.965 1.715 133.035 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 134.085 3.395 134.155 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 132.965 3.395 133.035 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 3.045 37.555 3.115 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 6.965 37.555 7.035 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 10.885 37.555 10.955 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 14.805 37.555 14.875 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 18.725 37.555 18.795 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 22.645 37.555 22.715 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 26.565 37.555 26.635 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 30.485 37.555 30.555 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 34.405 37.555 34.475 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 38.325 37.555 38.395 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 42.245 37.555 42.315 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 46.165 37.555 46.235 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 50.085 37.555 50.155 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 54.005 37.555 54.075 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 57.925 37.555 57.995 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 61.845 37.555 61.915 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 65.765 37.555 65.835 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 69.685 37.555 69.755 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 73.605 37.555 73.675 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 77.525 37.555 77.595 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 81.445 37.555 81.515 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 85.365 37.555 85.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 89.285 37.555 89.355 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 93.205 37.555 93.275 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 97.125 37.555 97.195 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 101.045 37.555 101.115 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 104.965 37.555 105.035 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 108.885 37.555 108.955 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 112.805 37.555 112.875 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 116.725 37.555 116.795 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 120.645 37.555 120.715 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 124.565 37.555 124.635 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 142.485 37.555 142.555 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 146.405 37.555 146.475 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 150.325 37.555 150.395 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 154.245 37.555 154.315 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 158.165 37.555 158.235 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 162.085 37.555 162.155 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 166.005 37.555 166.075 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 169.925 37.555 169.995 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 173.845 37.555 173.915 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 177.765 37.555 177.835 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 181.685 37.555 181.755 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 185.605 37.555 185.675 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 189.525 37.555 189.595 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 193.445 37.555 193.515 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 197.365 37.555 197.435 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 201.285 37.555 201.355 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 205.205 37.555 205.275 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 209.125 37.555 209.195 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 213.045 37.555 213.115 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 216.965 37.555 217.035 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 220.885 37.555 220.955 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 224.805 37.555 224.875 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 228.725 37.555 228.795 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 232.645 37.555 232.715 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 236.565 37.555 236.635 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 240.485 37.555 240.555 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 244.405 37.555 244.475 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 248.325 37.555 248.395 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 252.245 37.555 252.315 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 256.165 37.555 256.235 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 260.085 37.555 260.155 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 264.005 37.555 264.075 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 143.045 1.155 143.115 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 146.965 1.155 147.035 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 150.885 1.155 150.955 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 154.805 1.155 154.875 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 158.725 1.155 158.795 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 162.645 1.155 162.715 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 170.485 1.155 170.555 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.405 1.155 174.475 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.325 1.155 178.395 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.245 1.155 182.315 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.165 1.155 186.235 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.085 1.155 190.155 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.005 1.155 194.075 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 197.925 1.155 197.995 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 201.845 1.155 201.915 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 205.765 1.155 205.835 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 209.685 1.155 209.755 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 213.605 1.155 213.675 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 217.525 1.155 217.595 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 221.445 1.155 221.515 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.365 1.155 225.435 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.285 1.155 229.355 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.205 1.155 233.275 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.125 1.155 237.195 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.045 1.155 241.115 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 244.965 1.155 245.035 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 248.885 1.155 248.955 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 252.805 1.155 252.875 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 256.725 1.155 256.795 ;
        END
    END p271
    OBS
      LAYER via2 ;
        RECT  0 0 39.2 268.8 ;
      LAYER metal2 ;
        RECT  0 0 39.2 268.8 ;
      LAYER via1 ;
        RECT  0 0 39.2 268.8 ;
      LAYER metal1 ;
        RECT  0 0 39.2 268.8 ;
    END
END fake_macro_newblue1_o330459

MACRO fake_macro_newblue1_o330460
    CLASS BLOCK ;
    SIZE 53.76 BY 273.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 143.605 50.435 143.675 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 268.205 52.115 268.275 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 264.285 52.115 264.355 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 260.365 52.115 260.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 256.445 52.115 256.515 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 252.525 52.115 252.595 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 248.605 52.115 248.675 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 244.685 52.115 244.755 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 240.765 52.115 240.835 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 236.845 52.115 236.915 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 232.925 52.115 232.995 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 230.405 52.115 230.475 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 225.085 52.115 225.155 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 221.165 52.115 221.235 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 217.245 52.115 217.315 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 213.325 52.115 213.395 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 209.405 52.115 209.475 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 205.485 52.115 205.555 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 201.565 52.115 201.635 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 197.645 52.115 197.715 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 193.725 52.115 193.795 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 189.805 52.115 189.875 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 185.885 52.115 185.955 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 181.965 52.115 182.035 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 179.445 52.115 179.515 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 174.125 52.115 174.195 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 170.205 52.115 170.275 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 166.285 52.115 166.355 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 162.365 52.115 162.435 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 158.445 52.115 158.515 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 154.525 52.115 154.595 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 150.605 52.115 150.675 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 146.685 52.115 146.755 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 124.285 52.115 124.355 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 120.085 52.115 120.155 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 116.445 52.115 116.515 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 112.525 52.115 112.595 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 108.605 52.115 108.675 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 104.685 52.115 104.755 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 100.485 52.115 100.555 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 96.565 52.115 96.635 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 92.925 52.115 92.995 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 88.725 52.115 88.795 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 84.805 52.115 84.875 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 81.165 52.115 81.235 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 77.245 52.115 77.315 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 73.045 52.115 73.115 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 69.405 52.115 69.475 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 65.205 52.115 65.275 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 61.565 52.115 61.635 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 57.645 52.115 57.715 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 53.445 52.115 53.515 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 49.525 52.115 49.595 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 45.885 52.115 45.955 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 41.965 52.115 42.035 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 38.045 52.115 38.115 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 34.125 52.115 34.195 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 29.925 52.115 29.995 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 26.285 52.115 26.355 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 22.365 52.115 22.435 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 18.445 52.115 18.515 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 14.245 52.115 14.315 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 10.605 52.115 10.675 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 6.685 52.115 6.755 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 2.485 52.115 2.555 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.645 1.155 22.715 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.565 1.155 26.635 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.405 1.155 34.475 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 38.325 1.155 38.395 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.245 1.155 42.315 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.085 1.155 50.155 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 54.005 1.155 54.075 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.845 1.155 61.915 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.765 1.155 65.835 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.685 1.155 69.755 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.605 1.155 73.675 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 81.445 1.155 81.515 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 85.365 1.155 85.435 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.285 1.155 89.355 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 93.205 1.155 93.275 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.125 1.155 97.195 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 101.045 1.155 101.115 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.965 1.155 105.035 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.885 1.155 108.955 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.805 1.155 112.875 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.725 1.155 116.795 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.645 1.155 120.715 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.565 1.155 124.635 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 147.525 1.155 147.595 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.365 1.155 155.435 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.285 1.155 159.355 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 163.205 1.155 163.275 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 174.965 1.155 175.035 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 178.885 1.155 178.955 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 182.805 1.155 182.875 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 225.925 1.155 225.995 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 2.205 1.715 2.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 6.125 1.715 6.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 10.045 1.715 10.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 13.965 1.715 14.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 17.885 1.715 17.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 21.805 1.715 21.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 25.725 1.715 25.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 29.645 1.715 29.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 35.525 1.155 35.595 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 37.485 1.715 37.555 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 43.365 1.155 43.435 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 45.325 1.715 45.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 49.245 1.715 49.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 53.165 1.715 53.235 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 57.085 1.715 57.155 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 61.005 1.715 61.075 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 64.925 1.715 64.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 68.845 1.155 68.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 72.765 1.715 72.835 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 78.645 1.155 78.715 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 80.605 1.715 80.675 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 84.525 1.715 84.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 88.445 1.715 88.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 94.325 1.155 94.395 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 96.285 1.715 96.355 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 100.205 1.715 100.275 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 104.125 1.715 104.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 108.045 1.715 108.115 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 111.965 1.715 112.035 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 115.885 1.715 115.955 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 119.805 1.715 119.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 123.725 1.715 123.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 146.685 1.715 146.755 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 154.525 1.715 154.595 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 158.445 1.715 158.515 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 164.045 1.155 164.115 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 166.285 1.715 166.355 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.885 1.155 171.955 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 174.125 1.715 174.195 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 179.725 1.155 179.795 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 181.965 1.715 182.035 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 185.885 1.715 185.955 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 189.805 1.715 189.875 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 193.725 1.715 193.795 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 197.645 1.715 197.715 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 201.565 1.715 201.635 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 205.485 1.715 205.555 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 209.405 1.715 209.475 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.005 1.155 215.075 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 217.245 1.715 217.315 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 221.165 1.715 221.235 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 225.085 1.715 225.155 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 229.005 1.715 229.075 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 232.925 1.715 232.995 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 236.845 1.715 236.915 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 240.765 1.715 240.835 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 244.685 1.715 244.755 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 248.605 1.715 248.675 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 252.525 1.715 252.595 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 256.445 1.715 256.515 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 260.365 1.715 260.435 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 265.965 1.155 266.035 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 268.205 1.715 268.275 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 144.725 1.155 144.795 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 171.325 50.435 171.395 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 142.765 51.555 142.835 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 141.645 51.555 141.715 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 136.885 51.555 136.955 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 127.085 1.155 127.155 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.845 1.155 138.915 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 132.685 1.715 132.755 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 126.805 51.555 126.875 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 139.965 1.715 140.035 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.685 1.155 132.755 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 154.525 51.555 154.595 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 166.565 1.155 166.635 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 138.565 1.155 138.635 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.605 1.155 129.675 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 138.845 1.715 138.915 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 160.405 1.715 160.475 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 129.605 1.715 129.675 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 132.965 1.155 133.035 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 138.845 2.835 138.915 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.885 1.155 129.955 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.965 1.155 7.035 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.885 1.155 10.955 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.725 1.155 18.795 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 30.485 1.155 30.555 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 46.165 1.155 46.235 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.925 1.155 57.995 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 77.525 1.155 77.595 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 151.445 1.155 151.515 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 167.125 1.155 167.195 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.045 1.155 171.115 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 186.725 1.155 186.795 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 190.645 1.155 190.715 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 194.565 1.155 194.635 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 198.485 1.155 198.555 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.405 1.155 202.475 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.325 1.155 206.395 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 210.245 1.155 210.315 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 214.165 1.155 214.235 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 218.085 1.155 218.155 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 222.005 1.155 222.075 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 229.845 1.155 229.915 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 233.765 1.155 233.835 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 237.685 1.155 237.755 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 241.605 1.155 241.675 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 245.525 1.155 245.595 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 249.445 1.155 249.515 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.365 1.155 253.435 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.285 1.155 257.355 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 261.205 1.155 261.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 265.125 1.155 265.195 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 269.045 1.155 269.115 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 3.045 51.555 3.115 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 6.965 51.555 7.035 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 10.885 51.555 10.955 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 14.805 51.555 14.875 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 18.725 51.555 18.795 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 22.645 51.555 22.715 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 25.445 51.555 25.515 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 30.485 51.555 30.555 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 33.285 51.555 33.355 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 38.325 51.555 38.395 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 42.245 51.555 42.315 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 46.165 51.555 46.235 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 50.085 51.555 50.155 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 54.005 51.555 54.075 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 57.925 51.555 57.995 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 61.845 51.555 61.915 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 65.765 51.555 65.835 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 69.685 51.555 69.755 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 73.605 51.555 73.675 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 76.405 51.555 76.475 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 81.445 51.555 81.515 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 85.365 51.555 85.435 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 89.285 51.555 89.355 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 93.205 51.555 93.275 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 97.125 51.555 97.195 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 101.045 51.555 101.115 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 104.965 51.555 105.035 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 108.885 51.555 108.955 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 112.805 51.555 112.875 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 116.725 51.555 116.795 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 120.645 51.555 120.715 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 124.565 51.555 124.635 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 147.805 51.555 147.875 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 151.725 51.555 151.795 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 155.645 51.555 155.715 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 159.565 51.555 159.635 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 163.485 51.555 163.555 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 167.405 51.555 167.475 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 171.045 51.555 171.115 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 175.245 51.555 175.315 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 179.165 51.555 179.235 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 183.085 51.555 183.155 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 187.005 51.555 187.075 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 190.925 51.555 190.995 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 194.845 51.555 194.915 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 198.765 51.555 198.835 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 202.685 51.555 202.755 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 206.605 51.555 206.675 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 210.525 51.555 210.595 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 214.445 51.555 214.515 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 218.365 51.555 218.435 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 222.285 51.555 222.355 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 226.205 51.555 226.275 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 230.125 51.555 230.195 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 234.045 51.555 234.115 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 237.965 51.555 238.035 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 241.885 51.555 241.955 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 245.805 51.555 245.875 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 249.725 51.555 249.795 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 253.645 51.555 253.715 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 257.565 51.555 257.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 261.485 51.555 261.555 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 265.125 51.555 265.195 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 269.325 51.555 269.395 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.485 1.155 2.555 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 10.325 1.155 10.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.245 1.155 14.315 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 18.165 1.155 18.235 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.005 1.155 26.075 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 29.925 1.155 29.995 ;
        END
    END p285
    PIN p286
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 33.845 1.155 33.915 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 37.765 1.155 37.835 ;
        END
    END p287
    PIN p288
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 41.685 1.155 41.755 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 45.605 1.155 45.675 ;
        END
    END p289
    PIN p290
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 49.525 1.155 49.595 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 53.445 1.155 53.515 ;
        END
    END p291
    PIN p292
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 57.365 1.155 57.435 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 61.285 1.155 61.355 ;
        END
    END p293
    PIN p294
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 65.205 1.155 65.275 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 69.125 1.155 69.195 ;
        END
    END p295
    PIN p296
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.045 1.155 73.115 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 76.965 1.155 77.035 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 80.885 1.155 80.955 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 84.805 1.155 84.875 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 88.725 1.155 88.795 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 92.645 1.155 92.715 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 96.565 1.155 96.635 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 100.485 1.155 100.555 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 104.405 1.155 104.475 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 108.325 1.155 108.395 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 112.245 1.155 112.315 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 116.165 1.155 116.235 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 120.085 1.155 120.155 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 124.005 1.155 124.075 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 148.085 1.155 148.155 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 152.005 1.155 152.075 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 155.925 1.155 155.995 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 159.845 1.155 159.915 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 163.765 1.155 163.835 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 167.685 1.155 167.755 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 171.605 1.155 171.675 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 175.525 1.155 175.595 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 179.445 1.155 179.515 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 183.365 1.155 183.435 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 187.285 1.155 187.355 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 191.205 1.155 191.275 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 195.125 1.155 195.195 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 199.045 1.155 199.115 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 202.965 1.155 203.035 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 206.885 1.155 206.955 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 210.805 1.155 210.875 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 214.725 1.155 214.795 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 218.645 1.155 218.715 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 222.565 1.155 222.635 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 226.485 1.155 226.555 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 230.405 1.155 230.475 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 234.325 1.155 234.395 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 238.245 1.155 238.315 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 242.165 1.155 242.235 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 246.085 1.155 246.155 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 250.005 1.155 250.075 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 253.925 1.155 253.995 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 257.845 1.155 257.915 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 261.765 1.155 261.835 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 265.685 1.155 265.755 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 269.605 1.155 269.675 ;
        END
    END p341
    OBS
      LAYER via2 ;
        RECT  0 0 53.76 273.84 ;
      LAYER metal2 ;
        RECT  0 0 53.76 273.84 ;
      LAYER via1 ;
        RECT  0 0 53.76 273.84 ;
      LAYER metal1 ;
        RECT  0 0 53.76 273.84 ;
    END
END fake_macro_newblue1_o330460

MACRO fake_macro_newblue1_o330461
    CLASS BLOCK ;
    SIZE 132.16 BY 220.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 13.965 119.875 14.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 95.445 119.875 95.515 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  119.805 207.725 119.875 207.795 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 10.885 35.875 10.955 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 10.885 34.195 10.955 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 10.885 31.955 10.955 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 10.885 30.275 10.955 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 10.885 28.035 10.955 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.645 10.885 85.715 10.955 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 10.885 85.155 10.955 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 36.365 9.555 36.435 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 32.445 9.555 32.515 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 30.485 9.555 30.555 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 26.285 9.555 26.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 34.405 9.555 34.475 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 28.245 9.555 28.315 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 10.885 36.995 10.955 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  39.165 10.885 39.235 10.955 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 10.885 41.475 10.955 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 10.885 43.155 10.955 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 10.885 45.395 10.955 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 10.885 47.075 10.955 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 10.885 49.315 10.955 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 10.885 51.555 10.955 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 10.885 53.235 10.955 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  55.405 10.885 55.475 10.955 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 87.045 9.555 87.115 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 140.245 9.555 140.315 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 201.005 9.555 201.075 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 78.645 9.555 78.715 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 10.885 80.675 10.955 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 10.885 81.795 10.955 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 25.165 9.555 25.235 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 27.405 9.555 27.475 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 29.365 9.555 29.435 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 31.325 9.555 31.395 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 33.285 9.555 33.355 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 35.525 9.555 35.595 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 10.885 29.155 10.955 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 10.885 30.835 10.955 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 10.885 33.075 10.955 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 10.885 35.315 10.955 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  38.045 10.885 38.115 10.955 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.285 10.885 40.355 10.955 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 10.885 42.035 10.955 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 10.885 44.275 10.955 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  46.445 10.885 46.515 10.955 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 10.885 48.195 10.955 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 10.885 50.435 10.955 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 10.885 52.115 10.955 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 10.885 54.355 10.955 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 10.885 56.595 10.955 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 10.885 82.915 10.955 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 10.885 84.035 10.955 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 51.765 9.555 51.835 ;
        END
    END p54
    OBS
      LAYER via2 ;
        RECT  0 0 132.16 220.08 ;
      LAYER metal2 ;
        RECT  0 0 132.16 220.08 ;
      LAYER via1 ;
        RECT  0 0 132.16 220.08 ;
      LAYER metal1 ;
        RECT  0 0 132.16 220.08 ;
    END
END fake_macro_newblue1_o330461

MACRO fake_macro_newblue1_o330462
    CLASS BLOCK ;
    SIZE 132.16 BY 220.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 13.965 11.795 14.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 95.445 11.795 95.515 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 207.725 11.795 207.795 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 32.445 122.115 32.515 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 26.285 122.115 26.355 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 10.885 95.795 10.955 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 10.885 97.475 10.955 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.645 10.885 99.715 10.955 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 36.365 122.115 36.435 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 34.405 122.115 34.475 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 30.485 122.115 30.555 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 28.245 122.115 28.315 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.325 10.885 101.395 10.955 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 10.885 45.955 10.955 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  46.445 10.885 46.515 10.955 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 10.885 94.675 10.955 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  92.365 10.885 92.435 10.955 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.125 10.885 90.195 10.955 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  88.445 10.885 88.515 10.955 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 10.885 86.275 10.955 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  84.525 10.885 84.595 10.955 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 10.885 82.355 10.955 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 10.885 80.115 10.955 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.365 10.885 78.435 10.955 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 10.885 76.195 10.955 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.565 10.885 103.635 10.955 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 87.045 122.115 87.115 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 140.245 122.115 140.315 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 201.005 122.115 201.075 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 78.645 122.115 78.715 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 10.885 50.995 10.955 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 10.885 49.875 10.955 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 25.165 122.115 25.235 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 27.405 122.115 27.475 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 29.365 122.115 29.435 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 31.325 122.115 31.395 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 33.285 122.115 33.355 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 35.525 122.115 35.595 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 10.885 102.515 10.955 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  100.765 10.885 100.835 10.955 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 10.885 98.595 10.955 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 10.885 96.355 10.955 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 10.885 93.555 10.955 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 10.885 91.315 10.955 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.565 10.885 89.635 10.955 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 10.885 87.395 10.955 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 10.885 85.155 10.955 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 10.885 83.475 10.955 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.165 10.885 81.235 10.955 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 10.885 79.555 10.955 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.245 10.885 77.315 10.955 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 10.885 75.075 10.955 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 10.885 48.755 10.955 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.565 10.885 47.635 10.955 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  122.045 51.765 122.115 51.835 ;
        END
    END p54
    OBS
      LAYER via2 ;
        RECT  0 0 132.16 220.08 ;
      LAYER metal2 ;
        RECT  0 0 132.16 220.08 ;
      LAYER via1 ;
        RECT  0 0 132.16 220.08 ;
      LAYER metal1 ;
        RECT  0 0 132.16 220.08 ;
    END
END fake_macro_newblue1_o330462
END LIBRARY
