VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "|" ;

PROPERTYDEFINITIONS
END PROPERTYDEFINITIONS


MACRO fake_macro_adaptec1_o210904
    CLASS BLOCK ;
    SIZE 70 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.965 68.355 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.685 68.355 181.755 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 142.205 68.355 142.275 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.405 68.355 153.475 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 152.005 68.355 152.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.685 68.355 153.755 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 49.805 68.355 49.875 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 6.685 68.355 6.755 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 2.765 68.355 2.835 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 295.085 68.355 295.155 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 291.165 68.355 291.235 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 287.245 68.355 287.315 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 283.325 68.355 283.395 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 279.405 68.355 279.475 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 275.485 68.355 275.555 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 271.565 68.355 271.635 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 267.645 68.355 267.715 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 263.725 68.355 263.795 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 259.805 68.355 259.875 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 216.685 68.355 216.755 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 212.765 68.355 212.835 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 208.845 68.355 208.915 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 204.925 68.355 204.995 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 201.005 68.355 201.075 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 197.085 68.355 197.155 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 193.165 68.355 193.235 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 189.245 68.355 189.315 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 185.325 68.355 185.395 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.405 68.355 181.475 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 255.885 68.355 255.955 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 251.965 68.355 252.035 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 248.045 68.355 248.115 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 244.125 68.355 244.195 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 240.205 68.355 240.275 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 236.285 68.355 236.355 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 232.365 68.355 232.435 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 228.445 68.355 228.515 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 224.525 68.355 224.595 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 220.605 68.355 220.675 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 124.285 68.355 124.355 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 120.365 68.355 120.435 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 116.445 68.355 116.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 112.525 68.355 112.595 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 108.605 68.355 108.675 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 104.685 68.355 104.755 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 100.765 68.355 100.835 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 96.845 68.355 96.915 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 92.925 68.355 92.995 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 89.005 68.355 89.075 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 177.485 68.355 177.555 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 173.565 68.355 173.635 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.645 68.355 169.715 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 165.725 68.355 165.795 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 161.805 68.355 161.875 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 157.885 68.355 157.955 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 139.965 68.355 140.035 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 136.045 68.355 136.115 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 132.125 68.355 132.195 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 128.205 68.355 128.275 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 45.885 68.355 45.955 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 41.965 68.355 42.035 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 38.045 68.355 38.115 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 34.125 68.355 34.195 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 30.205 68.355 30.275 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 26.285 68.355 26.355 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 22.365 68.355 22.435 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 18.445 68.355 18.515 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 14.525 68.355 14.595 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 10.605 68.355 10.675 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 85.085 68.355 85.155 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 81.165 68.355 81.235 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 77.245 68.355 77.315 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 73.325 68.355 73.395 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.405 68.355 69.475 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 65.485 68.355 65.555 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 61.565 68.355 61.635 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 57.645 68.355 57.715 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 53.725 68.355 53.795 ;
        END
    END p377
    OBS
      LAYER via2 ;
        RECT  0 0 70 299.04 ;
      LAYER metal2 ;
        RECT  0 0 70 299.04 ;
      LAYER via1 ;
        RECT  0 0 70 299.04 ;
      LAYER metal1 ;
        RECT  0 0 70 299.04 ;
    END
END fake_macro_adaptec1_o210904

MACRO fake_macro_adaptec1_o210905
    CLASS BLOCK ;
    SIZE 70 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.965 68.355 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 142.205 68.355 142.275 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.925 68.355 169.995 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 152.005 68.355 152.075 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 154.245 68.915 154.315 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p285
    PIN p286
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p287
    PIN p288
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p289
    PIN p290
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p291
    PIN p292
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p293
    PIN p294
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p295
    PIN p296
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.685 68.355 153.755 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 6.685 68.355 6.755 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 2.765 68.355 2.835 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 216.685 68.355 216.755 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 212.765 68.355 212.835 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 208.845 68.355 208.915 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 204.925 68.355 204.995 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 201.005 68.355 201.075 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 197.085 68.355 197.155 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 193.165 68.355 193.235 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 189.245 68.355 189.315 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 185.325 68.355 185.395 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.405 68.355 181.475 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 255.885 68.355 255.955 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 251.965 68.355 252.035 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 248.045 68.355 248.115 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 244.125 68.355 244.195 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 240.205 68.355 240.275 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 236.285 68.355 236.355 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 232.365 68.355 232.435 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 228.445 68.355 228.515 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 224.525 68.355 224.595 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 220.605 68.355 220.675 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 124.285 68.355 124.355 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 120.365 68.355 120.435 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 116.445 68.355 116.515 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 112.525 68.355 112.595 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 108.605 68.355 108.675 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 104.685 68.355 104.755 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 100.765 68.355 100.835 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 96.845 68.355 96.915 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 92.925 68.355 92.995 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 89.005 68.355 89.075 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 177.485 68.355 177.555 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 173.565 68.355 173.635 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 295.085 68.355 295.155 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.645 68.355 169.715 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 291.165 68.355 291.235 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 165.725 68.355 165.795 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 287.245 68.355 287.315 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 161.805 68.355 161.875 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 283.325 68.355 283.395 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 157.885 68.355 157.955 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 279.405 68.355 279.475 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 139.965 68.355 140.035 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 275.485 68.355 275.555 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 136.045 68.355 136.115 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 271.565 68.355 271.635 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 132.125 68.355 132.195 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 267.645 68.355 267.715 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 128.205 68.355 128.275 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 263.725 68.355 263.795 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 259.805 68.355 259.875 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 45.885 68.355 45.955 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 41.965 68.355 42.035 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 38.045 68.355 38.115 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 34.125 68.355 34.195 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 30.205 68.355 30.275 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 26.285 68.355 26.355 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 22.365 68.355 22.435 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 18.445 68.355 18.515 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 14.525 68.355 14.595 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 10.605 68.355 10.675 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 85.085 68.355 85.155 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 81.165 68.355 81.235 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 77.245 68.355 77.315 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 73.325 68.355 73.395 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.405 68.355 69.475 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 65.485 68.355 65.555 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 61.565 68.355 61.635 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 57.645 68.355 57.715 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 53.725 68.355 53.795 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 49.805 68.355 49.875 ;
        END
    END p377
    OBS
      LAYER via2 ;
        RECT  0 0 70 299.04 ;
      LAYER metal2 ;
        RECT  0 0 70 299.04 ;
      LAYER via1 ;
        RECT  0 0 70 299.04 ;
      LAYER metal1 ;
        RECT  0 0 70 299.04 ;
    END
END fake_macro_adaptec1_o210905

MACRO fake_macro_adaptec1_o210906
    CLASS BLOCK ;
    SIZE 70 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.965 68.355 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.685 68.355 181.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 142.205 68.355 142.275 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.405 68.355 153.475 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 152.005 68.355 152.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.685 68.355 153.755 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 49.805 68.355 49.875 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 6.685 68.355 6.755 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 2.765 68.355 2.835 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 295.085 68.355 295.155 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 291.165 68.355 291.235 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 287.245 68.355 287.315 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 283.325 68.355 283.395 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 279.405 68.355 279.475 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 275.485 68.355 275.555 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 271.565 68.355 271.635 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 267.645 68.355 267.715 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 263.725 68.355 263.795 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 259.805 68.355 259.875 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 216.685 68.355 216.755 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 212.765 68.355 212.835 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 208.845 68.355 208.915 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 204.925 68.355 204.995 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 201.005 68.355 201.075 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 197.085 68.355 197.155 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 193.165 68.355 193.235 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 189.245 68.355 189.315 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 185.325 68.355 185.395 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.405 68.355 181.475 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 255.885 68.355 255.955 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 251.965 68.355 252.035 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 248.045 68.355 248.115 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 244.125 68.355 244.195 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 240.205 68.355 240.275 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 236.285 68.355 236.355 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 232.365 68.355 232.435 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 228.445 68.355 228.515 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 224.525 68.355 224.595 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 220.605 68.355 220.675 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 124.285 68.355 124.355 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 120.365 68.355 120.435 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 116.445 68.355 116.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 112.525 68.355 112.595 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 108.605 68.355 108.675 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 104.685 68.355 104.755 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 100.765 68.355 100.835 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 96.845 68.355 96.915 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 92.925 68.355 92.995 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 89.005 68.355 89.075 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 177.485 68.355 177.555 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 173.565 68.355 173.635 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.645 68.355 169.715 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 165.725 68.355 165.795 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 161.805 68.355 161.875 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 157.885 68.355 157.955 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 139.965 68.355 140.035 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 136.045 68.355 136.115 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 132.125 68.355 132.195 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 128.205 68.355 128.275 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 45.885 68.355 45.955 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 41.965 68.355 42.035 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 38.045 68.355 38.115 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 34.125 68.355 34.195 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 30.205 68.355 30.275 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 26.285 68.355 26.355 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 22.365 68.355 22.435 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 18.445 68.355 18.515 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 14.525 68.355 14.595 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 10.605 68.355 10.675 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 85.085 68.355 85.155 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 81.165 68.355 81.235 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 77.245 68.355 77.315 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 73.325 68.355 73.395 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.405 68.355 69.475 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 65.485 68.355 65.555 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 61.565 68.355 61.635 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 57.645 68.355 57.715 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 53.725 68.355 53.795 ;
        END
    END p377
    OBS
      LAYER via2 ;
        RECT  0 0 70 299.04 ;
      LAYER metal2 ;
        RECT  0 0 70 299.04 ;
      LAYER via1 ;
        RECT  0 0 70 299.04 ;
      LAYER metal1 ;
        RECT  0 0 70 299.04 ;
    END
END fake_macro_adaptec1_o210906

MACRO fake_macro_adaptec1_o210907
    CLASS BLOCK ;
    SIZE 70 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.965 68.355 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.685 68.355 181.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.685 68.355 153.755 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 142.205 68.355 142.275 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.405 68.355 153.475 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 152.005 68.355 152.075 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 6.685 68.355 6.755 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 2.765 68.355 2.835 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 216.685 68.355 216.755 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 212.765 68.355 212.835 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 208.845 68.355 208.915 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 204.925 68.355 204.995 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 201.005 68.355 201.075 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 197.085 68.355 197.155 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 193.165 68.355 193.235 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 189.245 68.355 189.315 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 185.325 68.355 185.395 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.405 68.355 181.475 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 255.885 68.355 255.955 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 251.965 68.355 252.035 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 248.045 68.355 248.115 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 244.125 68.355 244.195 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 240.205 68.355 240.275 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 236.285 68.355 236.355 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 232.365 68.355 232.435 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 228.445 68.355 228.515 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 224.525 68.355 224.595 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 220.605 68.355 220.675 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 124.285 68.355 124.355 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 120.365 68.355 120.435 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 116.445 68.355 116.515 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 112.525 68.355 112.595 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 108.605 68.355 108.675 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 104.685 68.355 104.755 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 100.765 68.355 100.835 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 96.845 68.355 96.915 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 92.925 68.355 92.995 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 89.005 68.355 89.075 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 177.485 68.355 177.555 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 173.565 68.355 173.635 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 295.085 68.355 295.155 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.645 68.355 169.715 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 291.165 68.355 291.235 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 165.725 68.355 165.795 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 287.245 68.355 287.315 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 161.805 68.355 161.875 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 283.325 68.355 283.395 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 157.885 68.355 157.955 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 279.405 68.355 279.475 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 139.965 68.355 140.035 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 275.485 68.355 275.555 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 136.045 68.355 136.115 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 271.565 68.355 271.635 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 132.125 68.355 132.195 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 267.645 68.355 267.715 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 128.205 68.355 128.275 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 263.725 68.355 263.795 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 259.805 68.355 259.875 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 45.885 68.355 45.955 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 41.965 68.355 42.035 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 38.045 68.355 38.115 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 34.125 68.355 34.195 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 30.205 68.355 30.275 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 26.285 68.355 26.355 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 22.365 68.355 22.435 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 18.445 68.355 18.515 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 14.525 68.355 14.595 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 10.605 68.355 10.675 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 85.085 68.355 85.155 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 81.165 68.355 81.235 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 77.245 68.355 77.315 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 73.325 68.355 73.395 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.405 68.355 69.475 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 65.485 68.355 65.555 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 61.565 68.355 61.635 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 57.645 68.355 57.715 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 53.725 68.355 53.795 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 49.805 68.355 49.875 ;
        END
    END p377
    OBS
      LAYER via2 ;
        RECT  0 0 70 299.04 ;
      LAYER metal2 ;
        RECT  0 0 70 299.04 ;
      LAYER via1 ;
        RECT  0 0 70 299.04 ;
      LAYER metal1 ;
        RECT  0 0 70 299.04 ;
    END
END fake_macro_adaptec1_o210907

MACRO fake_macro_adaptec1_o210908
    CLASS BLOCK ;
    SIZE 70 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.965 68.355 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.685 68.355 181.755 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 142.205 68.355 142.275 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.405 68.355 153.475 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 152.005 68.355 152.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.685 68.355 153.755 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 49.805 68.355 49.875 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 6.685 68.355 6.755 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 2.765 68.355 2.835 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 295.085 68.355 295.155 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 291.165 68.355 291.235 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 287.245 68.355 287.315 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 283.325 68.355 283.395 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 279.405 68.355 279.475 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 275.485 68.355 275.555 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 271.565 68.355 271.635 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 267.645 68.355 267.715 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 263.725 68.355 263.795 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 259.805 68.355 259.875 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 216.685 68.355 216.755 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 212.765 68.355 212.835 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 208.845 68.355 208.915 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 204.925 68.355 204.995 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 201.005 68.355 201.075 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 197.085 68.355 197.155 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 193.165 68.355 193.235 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 189.245 68.355 189.315 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 185.325 68.355 185.395 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.405 68.355 181.475 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 255.885 68.355 255.955 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 251.965 68.355 252.035 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 248.045 68.355 248.115 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 244.125 68.355 244.195 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 240.205 68.355 240.275 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 236.285 68.355 236.355 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 232.365 68.355 232.435 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 228.445 68.355 228.515 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 224.525 68.355 224.595 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 220.605 68.355 220.675 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 124.285 68.355 124.355 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 120.365 68.355 120.435 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 116.445 68.355 116.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 112.525 68.355 112.595 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 108.605 68.355 108.675 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 104.685 68.355 104.755 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 100.765 68.355 100.835 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 96.845 68.355 96.915 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 92.925 68.355 92.995 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 89.005 68.355 89.075 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 177.485 68.355 177.555 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 173.565 68.355 173.635 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.645 68.355 169.715 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 165.725 68.355 165.795 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 161.805 68.355 161.875 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 157.885 68.355 157.955 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 139.965 68.355 140.035 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 136.045 68.355 136.115 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 132.125 68.355 132.195 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 128.205 68.355 128.275 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 45.885 68.355 45.955 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 41.965 68.355 42.035 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 38.045 68.355 38.115 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 34.125 68.355 34.195 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 30.205 68.355 30.275 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 26.285 68.355 26.355 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 22.365 68.355 22.435 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 18.445 68.355 18.515 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 14.525 68.355 14.595 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 10.605 68.355 10.675 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 85.085 68.355 85.155 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 81.165 68.355 81.235 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 77.245 68.355 77.315 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 73.325 68.355 73.395 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.405 68.355 69.475 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 65.485 68.355 65.555 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 61.565 68.355 61.635 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 57.645 68.355 57.715 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 53.725 68.355 53.795 ;
        END
    END p377
    OBS
      LAYER via2 ;
        RECT  0 0 70 299.04 ;
      LAYER metal2 ;
        RECT  0 0 70 299.04 ;
      LAYER via1 ;
        RECT  0 0 70 299.04 ;
      LAYER metal1 ;
        RECT  0 0 70 299.04 ;
    END
END fake_macro_adaptec1_o210908

MACRO fake_macro_adaptec1_o210909
    CLASS BLOCK ;
    SIZE 70 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.965 68.355 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 142.205 68.355 142.275 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.925 68.355 169.995 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 152.005 68.355 152.075 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 154.245 68.915 154.315 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p285
    PIN p286
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p287
    PIN p288
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p289
    PIN p290
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p291
    PIN p292
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p293
    PIN p294
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p295
    PIN p296
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.685 68.355 153.755 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 6.685 68.355 6.755 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 2.765 68.355 2.835 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 216.685 68.355 216.755 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 212.765 68.355 212.835 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 208.845 68.355 208.915 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 204.925 68.355 204.995 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 201.005 68.355 201.075 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 197.085 68.355 197.155 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 193.165 68.355 193.235 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 189.245 68.355 189.315 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 185.325 68.355 185.395 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.405 68.355 181.475 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 255.885 68.355 255.955 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 251.965 68.355 252.035 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 248.045 68.355 248.115 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 244.125 68.355 244.195 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 240.205 68.355 240.275 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 236.285 68.355 236.355 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 232.365 68.355 232.435 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 228.445 68.355 228.515 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 224.525 68.355 224.595 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 220.605 68.355 220.675 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 124.285 68.355 124.355 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 120.365 68.355 120.435 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 116.445 68.355 116.515 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 112.525 68.355 112.595 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 108.605 68.355 108.675 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 104.685 68.355 104.755 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 100.765 68.355 100.835 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 96.845 68.355 96.915 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 92.925 68.355 92.995 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 89.005 68.355 89.075 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 177.485 68.355 177.555 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 173.565 68.355 173.635 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 295.085 68.355 295.155 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.645 68.355 169.715 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 291.165 68.355 291.235 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 165.725 68.355 165.795 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 287.245 68.355 287.315 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 161.805 68.355 161.875 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 283.325 68.355 283.395 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 157.885 68.355 157.955 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 279.405 68.355 279.475 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 139.965 68.355 140.035 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 275.485 68.355 275.555 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 136.045 68.355 136.115 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 271.565 68.355 271.635 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 132.125 68.355 132.195 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 267.645 68.355 267.715 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 128.205 68.355 128.275 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 263.725 68.355 263.795 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 259.805 68.355 259.875 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 45.885 68.355 45.955 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 41.965 68.355 42.035 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 38.045 68.355 38.115 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 34.125 68.355 34.195 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 30.205 68.355 30.275 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 26.285 68.355 26.355 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 22.365 68.355 22.435 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 18.445 68.355 18.515 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 14.525 68.355 14.595 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 10.605 68.355 10.675 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 85.085 68.355 85.155 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 81.165 68.355 81.235 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 77.245 68.355 77.315 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 73.325 68.355 73.395 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.405 68.355 69.475 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 65.485 68.355 65.555 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 61.565 68.355 61.635 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 57.645 68.355 57.715 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 53.725 68.355 53.795 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 49.805 68.355 49.875 ;
        END
    END p377
    OBS
      LAYER via2 ;
        RECT  0 0 70 299.04 ;
      LAYER metal2 ;
        RECT  0 0 70 299.04 ;
      LAYER via1 ;
        RECT  0 0 70 299.04 ;
      LAYER metal1 ;
        RECT  0 0 70 299.04 ;
    END
END fake_macro_adaptec1_o210909

MACRO fake_macro_adaptec1_o210910
    CLASS BLOCK ;
    SIZE 38.64 BY 146.16 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 75.565 36.995 75.635 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.045 0.595 143.115 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.605 0.595 129.675 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.685 0.595 125.755 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.925 0.595 113.995 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.405 0.595 90.475 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.485 0.595 86.555 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.685 0.595 62.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.405 0.595 27.475 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.925 0.595 78.995 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.045 0.595 80.115 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.845 0.595 82.915 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.965 0.595 84.035 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.765 0.595 86.835 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.885 0.595 87.955 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.685 0.595 90.755 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.805 0.595 91.875 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.605 0.595 94.675 ;
        END
    END p73
    PIN p74
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.725 0.595 95.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 98.525 0.595 98.595 ;
        END
    END p75
    PIN p76
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.645 0.595 99.715 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 102.445 0.595 102.515 ;
        END
    END p77
    PIN p78
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.565 0.595 103.635 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.365 0.595 106.435 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.285 0.595 110.355 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.405 0.595 111.475 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.205 0.595 114.275 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.325 0.595 115.395 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.125 0.595 118.195 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.245 0.595 119.315 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.045 0.595 122.115 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.165 0.595 123.235 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.965 0.595 126.035 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.085 0.595 127.155 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.885 0.595 129.955 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.005 0.595 131.075 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.805 0.595 133.875 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.925 0.595 134.995 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.725 0.595 137.795 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.845 0.595 138.915 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.645 0.595 141.715 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 73.605 36.995 73.675 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 71.085 0.595 71.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 71.085 1.715 71.155 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 71.085 2.835 71.155 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.205 0.595 142.275 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 63.805 36.995 63.875 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 91.525 36.995 91.595 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.965 0.595 70.035 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 69.965 1.715 70.035 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 69.965 2.835 70.035 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 75.845 37.555 75.915 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 75.285 36.995 75.355 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 79.485 0.595 79.555 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.405 0.595 83.475 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.325 0.595 87.395 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.245 0.595 91.315 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.165 0.595 95.235 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.085 0.595 99.155 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.005 0.595 103.075 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.925 0.595 106.995 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.845 0.595 110.915 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.765 0.595 114.835 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.685 0.595 118.755 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.605 0.595 122.675 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.525 0.595 126.595 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.445 0.595 130.515 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.365 0.595 134.435 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.285 0.595 138.355 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 45.885 36.995 45.955 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 41.965 36.995 42.035 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 38.045 36.995 38.115 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 34.125 36.995 34.195 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 30.205 36.995 30.275 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 26.285 36.995 26.355 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 22.365 36.995 22.435 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 18.445 36.995 18.515 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 14.525 36.995 14.595 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 10.605 36.995 10.675 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 99.085 36.995 99.155 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 95.165 36.995 95.235 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 91.245 36.995 91.315 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 87.325 36.995 87.395 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 83.405 36.995 83.475 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 79.485 36.995 79.555 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 61.565 36.995 61.635 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 57.645 36.995 57.715 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 53.725 36.995 53.795 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 49.805 36.995 49.875 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 138.285 36.995 138.355 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 134.365 36.995 134.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 130.445 36.995 130.515 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 126.525 36.995 126.595 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 122.605 36.995 122.675 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 118.685 36.995 118.755 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 114.765 36.995 114.835 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 110.845 36.995 110.915 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 106.925 36.995 106.995 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 103.005 36.995 103.075 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 6.685 36.995 6.755 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 2.765 36.995 2.835 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 142.205 36.995 142.275 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.485 0.595 107.555 ;
        END
    END p180
    OBS
      LAYER via2 ;
        RECT  0 0 38.64 146.16 ;
      LAYER metal2 ;
        RECT  0 0 38.64 146.16 ;
      LAYER via1 ;
        RECT  0 0 38.64 146.16 ;
      LAYER metal1 ;
        RECT  0 0 38.64 146.16 ;
    END
END fake_macro_adaptec1_o210910

MACRO fake_macro_adaptec1_o210911
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.925 21.315 169.995 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 154.245 21.875 154.315 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o210911

MACRO fake_macro_adaptec1_o210912
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.925 21.315 169.995 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 154.245 21.875 154.315 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o210912

MACRO fake_macro_adaptec1_o210913
    CLASS BLOCK ;
    SIZE 70 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.965 68.355 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.685 68.355 181.755 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 142.205 68.355 142.275 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.405 68.355 153.475 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 152.005 68.355 152.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.685 68.355 153.755 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 49.805 68.355 49.875 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 6.685 68.355 6.755 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 2.765 68.355 2.835 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 295.085 68.355 295.155 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 291.165 68.355 291.235 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 287.245 68.355 287.315 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 283.325 68.355 283.395 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 279.405 68.355 279.475 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 275.485 68.355 275.555 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 271.565 68.355 271.635 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 267.645 68.355 267.715 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 263.725 68.355 263.795 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 259.805 68.355 259.875 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 216.685 68.355 216.755 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 212.765 68.355 212.835 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 208.845 68.355 208.915 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 204.925 68.355 204.995 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 201.005 68.355 201.075 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 197.085 68.355 197.155 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 193.165 68.355 193.235 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 189.245 68.355 189.315 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 185.325 68.355 185.395 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.405 68.355 181.475 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 255.885 68.355 255.955 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 251.965 68.355 252.035 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 248.045 68.355 248.115 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 244.125 68.355 244.195 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 240.205 68.355 240.275 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 236.285 68.355 236.355 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 232.365 68.355 232.435 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 228.445 68.355 228.515 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 224.525 68.355 224.595 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 220.605 68.355 220.675 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 124.285 68.355 124.355 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 120.365 68.355 120.435 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 116.445 68.355 116.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 112.525 68.355 112.595 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 108.605 68.355 108.675 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 104.685 68.355 104.755 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 100.765 68.355 100.835 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 96.845 68.355 96.915 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 92.925 68.355 92.995 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 89.005 68.355 89.075 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 177.485 68.355 177.555 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 173.565 68.355 173.635 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.645 68.355 169.715 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 165.725 68.355 165.795 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 161.805 68.355 161.875 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 157.885 68.355 157.955 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 139.965 68.355 140.035 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 136.045 68.355 136.115 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 132.125 68.355 132.195 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 128.205 68.355 128.275 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 45.885 68.355 45.955 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 41.965 68.355 42.035 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 38.045 68.355 38.115 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 34.125 68.355 34.195 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 30.205 68.355 30.275 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 26.285 68.355 26.355 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 22.365 68.355 22.435 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 18.445 68.355 18.515 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 14.525 68.355 14.595 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 10.605 68.355 10.675 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 85.085 68.355 85.155 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 81.165 68.355 81.235 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 77.245 68.355 77.315 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 73.325 68.355 73.395 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.405 68.355 69.475 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 65.485 68.355 65.555 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 61.565 68.355 61.635 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 57.645 68.355 57.715 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 53.725 68.355 53.795 ;
        END
    END p377
    OBS
      LAYER via2 ;
        RECT  0 0 70 299.04 ;
      LAYER metal2 ;
        RECT  0 0 70 299.04 ;
      LAYER via1 ;
        RECT  0 0 70 299.04 ;
      LAYER metal1 ;
        RECT  0 0 70 299.04 ;
    END
END fake_macro_adaptec1_o210913

MACRO fake_macro_adaptec1_o210914
    CLASS BLOCK ;
    SIZE 70 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.965 68.355 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 153.685 68.355 153.755 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 142.205 68.355 142.275 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.925 68.355 169.995 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.525 2.275 147.595 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 152.005 68.355 152.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 150.605 1.715 150.675 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 154.245 68.915 154.315 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 6.685 68.355 6.755 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 2.765 68.355 2.835 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 216.685 68.355 216.755 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 212.765 68.355 212.835 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 208.845 68.355 208.915 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 204.925 68.355 204.995 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 201.005 68.355 201.075 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 197.085 68.355 197.155 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 193.165 68.355 193.235 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 189.245 68.355 189.315 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 185.325 68.355 185.395 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 181.405 68.355 181.475 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 255.885 68.355 255.955 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 251.965 68.355 252.035 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 248.045 68.355 248.115 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 244.125 68.355 244.195 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 240.205 68.355 240.275 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 236.285 68.355 236.355 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 232.365 68.355 232.435 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 228.445 68.355 228.515 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 224.525 68.355 224.595 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 220.605 68.355 220.675 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 124.285 68.355 124.355 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 120.365 68.355 120.435 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 116.445 68.355 116.515 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 112.525 68.355 112.595 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 108.605 68.355 108.675 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 104.685 68.355 104.755 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 100.765 68.355 100.835 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 96.845 68.355 96.915 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 92.925 68.355 92.995 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 89.005 68.355 89.075 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 177.485 68.355 177.555 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 173.565 68.355 173.635 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 295.085 68.355 295.155 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 169.645 68.355 169.715 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 291.165 68.355 291.235 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 165.725 68.355 165.795 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 287.245 68.355 287.315 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 161.805 68.355 161.875 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 283.325 68.355 283.395 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 157.885 68.355 157.955 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 279.405 68.355 279.475 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 139.965 68.355 140.035 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 275.485 68.355 275.555 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 136.045 68.355 136.115 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 271.565 68.355 271.635 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 132.125 68.355 132.195 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 267.645 68.355 267.715 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 128.205 68.355 128.275 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 263.725 68.355 263.795 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 259.805 68.355 259.875 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 45.885 68.355 45.955 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 41.965 68.355 42.035 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 38.045 68.355 38.115 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 34.125 68.355 34.195 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 30.205 68.355 30.275 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 26.285 68.355 26.355 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 22.365 68.355 22.435 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 18.445 68.355 18.515 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 14.525 68.355 14.595 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 10.605 68.355 10.675 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 85.085 68.355 85.155 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 81.165 68.355 81.235 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 77.245 68.355 77.315 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 73.325 68.355 73.395 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 69.405 68.355 69.475 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 65.485 68.355 65.555 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 61.565 68.355 61.635 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 57.645 68.355 57.715 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 53.725 68.355 53.795 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 49.805 68.355 49.875 ;
        END
    END p377
    OBS
      LAYER via2 ;
        RECT  0 0 70 299.04 ;
      LAYER metal2 ;
        RECT  0 0 70 299.04 ;
      LAYER via1 ;
        RECT  0 0 70 299.04 ;
      LAYER metal1 ;
        RECT  0 0 70 299.04 ;
    END
END fake_macro_adaptec1_o210914

MACRO fake_macro_adaptec1_o210915
    CLASS BLOCK ;
    SIZE 168.84 BY 399.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 11.165 2.835 11.235 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 21.525 2.835 21.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 23.765 3.395 23.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 23.765 2.835 23.835 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 26.005 3.395 26.075 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 26.005 2.835 26.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 28.245 3.395 28.315 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 28.245 2.835 28.315 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 30.485 3.395 30.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 30.485 2.835 30.555 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 17.045 3.395 17.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 17.045 2.835 17.115 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 19.285 3.395 19.355 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 19.285 2.835 19.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.525 3.395 21.595 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 4.725 11.795 4.795 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 4.725 14.595 4.795 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 4.725 14.035 4.795 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 4.725 15.715 4.795 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.285 1.715 12.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 5.845 5.075 5.915 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 5.845 7.315 5.915 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 1.085 6.195 1.155 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 1.085 11.235 1.155 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 32.445 11.795 32.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 1.085 22.435 1.155 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 1.085 26.355 1.155 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 1.085 29.715 1.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 1.085 33.635 1.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 1.085 41.475 1.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 1.085 44.835 1.155 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 1.085 48.755 1.155 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 1.085 52.115 1.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.085 57.155 1.155 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 1.085 60.515 1.155 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 1.085 64.435 1.155 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 1.085 67.795 1.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 1.085 75.635 1.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 1.085 79.555 1.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 1.085 82.915 1.155 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 1.085 86.835 1.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 1.085 91.315 1.155 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 1.085 95.235 1.155 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 1.085 98.595 1.155 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 1.085 102.515 1.155 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.285 1.085 110.355 1.155 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.645 1.085 113.715 1.155 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.565 1.085 117.635 1.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 1.085 120.995 1.155 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 1.085 126.035 1.155 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.325 1.085 129.395 1.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 1.085 133.315 1.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.605 1.085 136.675 1.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  144.445 1.085 144.515 1.155 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.365 1.085 148.435 1.155 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.725 1.085 151.795 1.155 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.645 1.085 155.715 1.155 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 49.245 3.395 49.315 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.245 3.395 21.315 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 19.565 3.955 19.635 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 19.005 3.955 19.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.765 3.955 30.835 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.205 3.955 30.275 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 28.525 3.955 28.595 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 27.965 3.955 28.035 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 26.285 3.955 26.355 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 25.725 3.955 25.795 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 24.045 3.955 24.115 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 23.485 3.955 23.555 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 11.165 3.395 11.235 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 4.725 12.915 4.795 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.125 1.085 160.195 1.155 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 12.285 12.355 12.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 1.085 48.195 1.155 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 1.085 44.275 1.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.845 1.085 40.915 1.155 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 1.085 33.075 1.155 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 1.085 29.155 1.155 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 1.085 25.795 1.155 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 1.085 21.875 1.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  128.765 1.085 128.835 1.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 1.085 90.755 1.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.085 51.555 1.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.885 1.085 101.955 1.155 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.965 1.085 98.035 1.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 1.085 94.675 1.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 1.085 86.275 1.155 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 1.085 82.355 1.155 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 1.085 78.995 1.155 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 1.085 75.075 1.155 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 1.085 67.235 1.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 1.085 63.875 1.155 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.885 1.085 59.955 1.155 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 1.085 56.595 1.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 1.085 159.635 1.155 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.085 1.085 155.155 1.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.165 1.085 151.235 1.155 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.805 1.085 147.875 1.155 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  143.885 1.085 143.955 1.155 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 1.085 136.115 1.155 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.685 1.085 132.755 1.155 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.405 1.085 125.475 1.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 1.085 120.435 1.155 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 1.085 117.075 1.155 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.085 1.085 113.155 1.155 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  109.725 1.085 109.795 1.155 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.685 17.325 160.755 17.395 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  156.205 17.325 156.275 17.395 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.285 17.325 152.355 17.395 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.925 17.325 148.995 17.395 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.005 17.325 145.075 17.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.165 17.325 137.235 17.395 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.805 17.325 133.875 17.395 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.885 17.325 129.955 17.395 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  126.525 17.325 126.595 17.395 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 17.325 121.555 17.395 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.125 17.325 118.195 17.395 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.565 1.715 12.635 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.205 17.325 114.275 17.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.845 17.325 110.915 17.395 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 17.325 103.075 17.395 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 17.325 99.155 17.395 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 17.325 95.795 17.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 17.325 91.875 17.395 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 17.325 87.395 17.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 17.325 83.475 17.395 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 17.325 80.115 17.395 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 17.325 76.195 17.395 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 17.325 68.355 17.395 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 17.325 64.995 17.395 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 17.325 61.075 17.395 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 17.325 57.715 17.395 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 17.325 52.675 17.395 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 17.325 49.315 17.395 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 17.325 45.395 17.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 17.325 42.035 17.395 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 17.325 34.195 17.395 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 17.325 30.275 17.395 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 17.325 26.915 17.395 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 17.325 22.995 17.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 19.565 10.115 19.635 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.845 1.715 12.915 ;
        END
    END p141
    OBS
      LAYER via2 ;
        RECT  0 0 168.84 399.84 ;
      LAYER metal2 ;
        RECT  0 0 168.84 399.84 ;
      LAYER via1 ;
        RECT  0 0 168.84 399.84 ;
      LAYER metal1 ;
        RECT  0 0 168.84 399.84 ;
    END
END fake_macro_adaptec1_o210915

MACRO fake_macro_adaptec1_o210916
    CLASS BLOCK ;
    SIZE 168.84 BY 399.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 11.165 2.835 11.235 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 21.525 2.835 21.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 23.765 3.395 23.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 23.765 2.835 23.835 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 26.005 3.395 26.075 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 26.005 2.835 26.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 28.245 3.395 28.315 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 28.245 2.835 28.315 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 30.485 3.395 30.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 30.485 2.835 30.555 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 17.045 3.395 17.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 17.045 2.835 17.115 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 19.285 3.395 19.355 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 19.285 2.835 19.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.525 3.395 21.595 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 4.725 11.795 4.795 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 4.725 14.595 4.795 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 4.725 14.035 4.795 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 4.725 15.715 4.795 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.285 1.715 12.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 5.845 5.075 5.915 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 5.845 7.315 5.915 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 1.085 6.195 1.155 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 1.085 11.235 1.155 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 32.445 11.795 32.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 49.245 3.395 49.315 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.245 3.395 21.315 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 19.565 3.955 19.635 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 19.005 3.955 19.075 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.765 3.955 30.835 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.205 3.955 30.275 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 28.525 3.955 28.595 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 27.965 3.955 28.035 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 26.285 3.955 26.355 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 25.725 3.955 25.795 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 24.045 3.955 24.115 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 23.485 3.955 23.555 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 12.285 12.355 12.355 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 1.085 22.435 1.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 1.085 26.355 1.155 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 1.085 29.715 1.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 1.085 33.635 1.155 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 1.085 41.475 1.155 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 1.085 44.835 1.155 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 1.085 48.755 1.155 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 1.085 52.115 1.155 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.085 57.155 1.155 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 1.085 60.515 1.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 1.085 64.435 1.155 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 1.085 67.795 1.155 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 1.085 75.635 1.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 1.085 79.555 1.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 1.085 82.915 1.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 1.085 86.835 1.155 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 1.085 91.315 1.155 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 1.085 95.235 1.155 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 1.085 98.595 1.155 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 1.085 102.515 1.155 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.285 1.085 110.355 1.155 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.645 1.085 113.715 1.155 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.565 1.085 117.635 1.155 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 1.085 120.995 1.155 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 1.085 126.035 1.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.325 1.085 129.395 1.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 1.085 133.315 1.155 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.605 1.085 136.675 1.155 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  144.445 1.085 144.515 1.155 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.365 1.085 148.435 1.155 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.725 1.085 151.795 1.155 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.645 1.085 155.715 1.155 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 11.165 3.395 11.235 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 4.725 12.915 4.795 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.125 1.085 160.195 1.155 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 1.085 33.075 1.155 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 1.085 29.155 1.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 1.085 21.875 1.155 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  143.885 1.085 143.955 1.155 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.885 1.085 101.955 1.155 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 1.085 63.875 1.155 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 1.085 25.795 1.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.965 1.085 98.035 1.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 1.085 94.675 1.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 1.085 90.755 1.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 1.085 86.275 1.155 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 1.085 82.355 1.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 1.085 78.995 1.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 1.085 75.075 1.155 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 1.085 67.235 1.155 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.885 1.085 59.955 1.155 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 1.085 56.595 1.155 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.085 51.555 1.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 1.085 48.195 1.155 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 1.085 44.275 1.155 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.845 1.085 40.915 1.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 1.085 159.635 1.155 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.085 1.085 155.155 1.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.165 1.085 151.235 1.155 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.805 1.085 147.875 1.155 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 1.085 136.115 1.155 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.685 1.085 132.755 1.155 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  128.765 1.085 128.835 1.155 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.405 1.085 125.475 1.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 1.085 120.435 1.155 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 1.085 117.075 1.155 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.085 1.085 113.155 1.155 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  109.725 1.085 109.795 1.155 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.845 1.715 12.915 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.685 17.325 160.755 17.395 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.565 1.715 12.635 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  156.205 17.325 156.275 17.395 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.285 17.325 152.355 17.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.925 17.325 148.995 17.395 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.005 17.325 145.075 17.395 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.165 17.325 137.235 17.395 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.805 17.325 133.875 17.395 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.885 17.325 129.955 17.395 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  126.525 17.325 126.595 17.395 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 17.325 121.555 17.395 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.125 17.325 118.195 17.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.205 17.325 114.275 17.395 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.845 17.325 110.915 17.395 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 17.325 103.075 17.395 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 17.325 99.155 17.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 17.325 95.795 17.395 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 17.325 91.875 17.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 17.325 87.395 17.395 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 17.325 83.475 17.395 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 17.325 80.115 17.395 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 17.325 76.195 17.395 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 17.325 68.355 17.395 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 17.325 64.995 17.395 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 17.325 61.075 17.395 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 17.325 57.715 17.395 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 17.325 52.675 17.395 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 17.325 49.315 17.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 17.325 45.395 17.395 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 17.325 42.035 17.395 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 17.325 34.195 17.395 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 17.325 30.275 17.395 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 17.325 26.915 17.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 17.325 22.995 17.395 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 19.565 10.115 19.635 ;
        END
    END p141
    OBS
      LAYER via2 ;
        RECT  0 0 168.84 399.84 ;
      LAYER metal2 ;
        RECT  0 0 168.84 399.84 ;
      LAYER via1 ;
        RECT  0 0 168.84 399.84 ;
      LAYER metal1 ;
        RECT  0 0 168.84 399.84 ;
    END
END fake_macro_adaptec1_o210916

MACRO fake_macro_adaptec1_o210917
    CLASS BLOCK ;
    SIZE 168.84 BY 399.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 11.165 2.835 11.235 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 21.525 2.835 21.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 23.765 3.395 23.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 23.765 2.835 23.835 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 26.005 3.395 26.075 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 26.005 2.835 26.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 28.245 3.395 28.315 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 28.245 2.835 28.315 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 30.485 3.395 30.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 30.485 2.835 30.555 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 17.045 3.395 17.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 17.045 2.835 17.115 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 19.285 3.395 19.355 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 19.285 2.835 19.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.525 3.395 21.595 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 4.725 11.795 4.795 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 4.725 14.595 4.795 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 4.725 14.035 4.795 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 4.725 15.715 4.795 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.285 1.715 12.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 5.845 5.075 5.915 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 5.845 7.315 5.915 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 1.085 6.195 1.155 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 32.445 11.795 32.515 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 1.085 22.435 1.155 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 1.085 26.355 1.155 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 1.085 29.715 1.155 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 1.085 33.635 1.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 1.085 41.475 1.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 1.085 44.835 1.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 1.085 48.755 1.155 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 1.085 52.115 1.155 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.085 57.155 1.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 1.085 60.515 1.155 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 1.085 64.435 1.155 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 1.085 67.795 1.155 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 1.085 75.635 1.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 1.085 79.555 1.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 1.085 82.915 1.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 1.085 86.835 1.155 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 1.085 91.315 1.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 1.085 95.235 1.155 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 1.085 98.595 1.155 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 1.085 102.515 1.155 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.285 1.085 110.355 1.155 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.645 1.085 113.715 1.155 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.565 1.085 117.635 1.155 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 1.085 120.995 1.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 1.085 126.035 1.155 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.325 1.085 129.395 1.155 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 1.085 133.315 1.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.605 1.085 136.675 1.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  144.445 1.085 144.515 1.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.365 1.085 148.435 1.155 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.725 1.085 151.795 1.155 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.645 1.085 155.715 1.155 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 49.245 3.395 49.315 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.245 3.395 21.315 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 19.565 3.955 19.635 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 19.005 3.955 19.075 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.765 3.955 30.835 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.205 3.955 30.275 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 28.525 3.955 28.595 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 27.965 3.955 28.035 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 26.285 3.955 26.355 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 25.725 3.955 25.795 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 24.045 3.955 24.115 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 23.485 3.955 23.555 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 11.165 3.395 11.235 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.125 1.085 160.195 1.155 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 12.285 12.355 12.355 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 1.085 11.235 1.155 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 4.725 12.915 4.795 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 1.085 67.235 1.155 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 1.085 63.875 1.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.885 1.085 59.955 1.155 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 1.085 56.595 1.155 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.085 51.555 1.155 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 1.085 48.195 1.155 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 1.085 44.275 1.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 1.085 33.075 1.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 1.085 29.155 1.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 1.085 25.795 1.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 1.085 21.875 1.155 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 1.085 117.075 1.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.085 1.085 113.155 1.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 1.085 78.995 1.155 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.845 1.085 40.915 1.155 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 1.085 120.435 1.155 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  109.725 1.085 109.795 1.155 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.885 1.085 101.955 1.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.965 1.085 98.035 1.155 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 1.085 94.675 1.155 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 1.085 90.755 1.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 1.085 86.275 1.155 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 1.085 82.355 1.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 1.085 75.075 1.155 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 1.085 159.635 1.155 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.085 1.085 155.155 1.155 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.165 1.085 151.235 1.155 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.805 1.085 147.875 1.155 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  143.885 1.085 143.955 1.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 1.085 136.115 1.155 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.685 1.085 132.755 1.155 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  128.765 1.085 128.835 1.155 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.405 1.085 125.475 1.155 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.565 1.715 12.635 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.845 1.715 12.915 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.685 17.325 160.755 17.395 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  156.205 17.325 156.275 17.395 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.285 17.325 152.355 17.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.925 17.325 148.995 17.395 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.005 17.325 145.075 17.395 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.165 17.325 137.235 17.395 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.805 17.325 133.875 17.395 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.885 17.325 129.955 17.395 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  126.525 17.325 126.595 17.395 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 17.325 121.555 17.395 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.125 17.325 118.195 17.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.205 17.325 114.275 17.395 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.845 17.325 110.915 17.395 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 17.325 103.075 17.395 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 17.325 99.155 17.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 17.325 95.795 17.395 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 17.325 91.875 17.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 17.325 87.395 17.395 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 17.325 83.475 17.395 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 17.325 80.115 17.395 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 17.325 76.195 17.395 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 17.325 68.355 17.395 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 17.325 64.995 17.395 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 17.325 61.075 17.395 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 17.325 57.715 17.395 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 17.325 52.675 17.395 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 17.325 49.315 17.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 17.325 45.395 17.395 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 17.325 42.035 17.395 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 17.325 34.195 17.395 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 17.325 30.275 17.395 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 17.325 26.915 17.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 17.325 22.995 17.395 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 19.565 10.115 19.635 ;
        END
    END p141
    OBS
      LAYER via2 ;
        RECT  0 0 168.84 399.84 ;
      LAYER metal2 ;
        RECT  0 0 168.84 399.84 ;
      LAYER via1 ;
        RECT  0 0 168.84 399.84 ;
      LAYER metal1 ;
        RECT  0 0 168.84 399.84 ;
    END
END fake_macro_adaptec1_o210917

MACRO fake_macro_adaptec1_o210918
    CLASS BLOCK ;
    SIZE 168.84 BY 399.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.525 3.395 21.595 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 49.245 3.395 49.315 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 19.285 3.395 19.355 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.245 3.395 21.315 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 30.485 3.395 30.555 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.765 3.955 30.835 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 28.245 3.395 28.315 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 28.525 3.955 28.595 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 26.005 3.395 26.075 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 26.285 3.955 26.355 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 23.765 3.395 23.835 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 24.045 3.955 24.115 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 1.085 22.435 1.155 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 1.085 26.355 1.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 1.085 29.715 1.155 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 1.085 33.635 1.155 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 1.085 41.475 1.155 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 1.085 44.835 1.155 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 1.085 48.755 1.155 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 1.085 52.115 1.155 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.085 57.155 1.155 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 1.085 60.515 1.155 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 1.085 64.435 1.155 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 1.085 67.795 1.155 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 1.085 75.635 1.155 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 1.085 79.555 1.155 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 1.085 82.915 1.155 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 1.085 86.835 1.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 1.085 91.315 1.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 1.085 95.235 1.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 1.085 98.595 1.155 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 1.085 102.515 1.155 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.285 1.085 110.355 1.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.645 1.085 113.715 1.155 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.565 1.085 117.635 1.155 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.925 1.085 120.995 1.155 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 1.085 126.035 1.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.325 1.085 129.395 1.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.245 1.085 133.315 1.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.605 1.085 136.675 1.155 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  144.445 1.085 144.515 1.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.365 1.085 148.435 1.155 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.725 1.085 151.795 1.155 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.645 1.085 155.715 1.155 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 11.165 3.395 11.235 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.125 1.085 160.195 1.155 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 12.285 12.355 12.355 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 1.085 11.235 1.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 11.165 2.835 11.235 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 21.525 2.835 21.595 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 23.485 3.955 23.555 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 23.765 2.835 23.835 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 25.725 3.955 25.795 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 26.005 2.835 26.075 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 27.965 3.955 28.035 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 28.245 2.835 28.315 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.205 3.955 30.275 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 30.485 2.835 30.555 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 17.045 3.395 17.115 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 17.045 2.835 17.115 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 19.565 3.955 19.635 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 19.285 2.835 19.355 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 21.805 3.955 21.875 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 4.725 11.795 4.795 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 4.725 14.595 4.795 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 4.725 14.035 4.795 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 4.725 15.715 4.795 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.285 1.715 12.355 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 5.845 5.075 5.915 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 5.845 7.315 5.915 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 1.085 6.195 1.155 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 32.445 11.795 32.515 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 4.725 12.915 4.795 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 1.085 33.075 1.155 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 1.085 29.155 1.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 1.085 25.795 1.155 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 1.085 21.875 1.155 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 1.085 67.235 1.155 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 1.085 63.875 1.155 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.885 1.085 59.955 1.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 1.085 56.595 1.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.085 51.555 1.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 1.085 48.195 1.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 1.085 44.275 1.155 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.845 1.085 40.915 1.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  101.885 1.085 101.955 1.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.965 1.085 98.035 1.155 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 1.085 94.675 1.155 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 1.085 90.755 1.155 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 1.085 86.275 1.155 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 1.085 82.355 1.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 1.085 78.995 1.155 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 1.085 75.075 1.155 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 1.085 136.115 1.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  132.685 1.085 132.755 1.155 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  128.765 1.085 128.835 1.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.405 1.085 125.475 1.155 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  120.365 1.085 120.435 1.155 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  117.005 1.085 117.075 1.155 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  113.085 1.085 113.155 1.155 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  109.725 1.085 109.795 1.155 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  159.565 1.085 159.635 1.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  155.085 1.085 155.155 1.155 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  151.165 1.085 151.235 1.155 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  147.805 1.085 147.875 1.155 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  143.885 1.085 143.955 1.155 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 19.565 10.115 19.635 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  160.685 17.325 160.755 17.395 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.845 1.715 12.915 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  156.205 17.325 156.275 17.395 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  152.285 17.325 152.355 17.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  148.925 17.325 148.995 17.395 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  145.005 17.325 145.075 17.395 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  137.165 17.325 137.235 17.395 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  133.805 17.325 133.875 17.395 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  129.885 17.325 129.955 17.395 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  126.525 17.325 126.595 17.395 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  121.485 17.325 121.555 17.395 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  118.125 17.325 118.195 17.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  114.205 17.325 114.275 17.395 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  110.845 17.325 110.915 17.395 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 17.325 103.075 17.395 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 17.325 99.155 17.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 17.325 95.795 17.395 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 17.325 91.875 17.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 17.325 87.395 17.395 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 17.325 83.475 17.395 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 17.325 80.115 17.395 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 17.325 76.195 17.395 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 17.325 68.355 17.395 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 17.325 64.995 17.395 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 17.325 61.075 17.395 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 17.325 57.715 17.395 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 17.325 52.675 17.395 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 17.325 49.315 17.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 17.325 45.395 17.395 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 17.325 42.035 17.395 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 17.325 34.195 17.395 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 17.325 30.275 17.395 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 17.325 26.915 17.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 17.325 22.995 17.395 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.565 1.715 12.635 ;
        END
    END p141
    OBS
      LAYER via2 ;
        RECT  0 0 168.84 399.84 ;
      LAYER metal2 ;
        RECT  0 0 168.84 399.84 ;
      LAYER via1 ;
        RECT  0 0 168.84 399.84 ;
      LAYER metal1 ;
        RECT  0 0 168.84 399.84 ;
    END
END fake_macro_adaptec1_o210918

MACRO fake_macro_adaptec1_o210919
    CLASS BLOCK ;
    SIZE 11.2 BY 146.16 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 63.805 9.555 63.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.205 0.595 142.275 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.285 0.595 138.355 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.365 0.595 134.435 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.445 0.595 130.515 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.525 0.595 126.595 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.605 0.595 122.675 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.685 0.595 118.755 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.765 0.595 114.835 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.845 0.595 110.915 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.925 0.595 106.995 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.005 0.595 103.075 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.085 0.595 99.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.165 0.595 95.235 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.245 0.595 91.315 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.325 0.595 87.395 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.405 0.595 83.475 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 79.485 0.595 79.555 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 75.565 9.555 75.635 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.045 0.595 143.115 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.605 0.595 129.675 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.765 0.595 121.835 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.925 0.595 113.995 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.325 0.595 94.395 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.485 0.595 86.555 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.685 0.595 62.755 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.405 0.595 27.475 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 91.525 9.555 91.595 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 75.845 10.115 75.915 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p74
    PIN p75
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.925 0.595 78.995 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.045 0.595 80.115 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.845 0.595 82.915 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.965 0.595 84.035 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.765 0.595 86.835 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.885 0.595 87.955 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.685 0.595 90.755 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.805 0.595 91.875 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.605 0.595 94.675 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.725 0.595 95.795 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 98.525 0.595 98.595 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.645 0.595 99.715 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 102.445 0.595 102.515 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.565 0.595 103.635 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.365 0.595 106.435 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.485 0.595 107.555 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.285 0.595 110.355 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.405 0.595 111.475 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.205 0.595 114.275 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.325 0.595 115.395 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.125 0.595 118.195 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.245 0.595 119.315 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.045 0.595 122.115 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.165 0.595 123.235 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.965 0.595 126.035 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.085 0.595 127.155 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.885 0.595 129.955 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.005 0.595 131.075 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.805 0.595 133.875 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.925 0.595 134.995 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.725 0.595 137.795 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.845 0.595 138.915 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.645 0.595 141.715 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 73.605 9.555 73.675 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 75.285 9.555 75.355 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 142.205 9.555 142.275 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.285 9.555 138.355 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 134.365 9.555 134.435 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 126.525 9.555 126.595 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 122.605 9.555 122.675 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.605 9.555 10.675 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 118.685 9.555 118.755 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 6.685 9.555 6.755 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 114.765 9.555 114.835 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.765 9.555 2.835 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 110.845 9.555 110.915 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 106.925 9.555 106.995 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 49.805 9.555 49.875 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 45.885 9.555 45.955 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 38.045 9.555 38.115 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 34.125 9.555 34.195 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 30.205 9.555 30.275 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 26.285 9.555 26.355 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 22.365 9.555 22.435 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 18.445 9.555 18.515 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 14.525 9.555 14.595 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 103.005 9.555 103.075 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 99.085 9.555 99.155 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 95.165 9.555 95.235 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 91.245 9.555 91.315 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 87.325 9.555 87.395 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 83.405 9.555 83.475 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 79.485 9.555 79.555 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 61.565 9.555 61.635 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 57.645 9.555 57.715 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 53.725 9.555 53.795 ;
        END
    END p174
    OBS
      LAYER via2 ;
        RECT  0 0 11.2 146.16 ;
      LAYER metal2 ;
        RECT  0 0 11.2 146.16 ;
      LAYER via1 ;
        RECT  0 0 11.2 146.16 ;
      LAYER metal1 ;
        RECT  0 0 11.2 146.16 ;
    END
END fake_macro_adaptec1_o210919

MACRO fake_macro_adaptec1_o210920
    CLASS BLOCK ;
    SIZE 38.64 BY 307.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 152.285 0.595 152.355 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 146.125 36.995 146.195 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 173.845 36.995 173.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 147.245 0.595 147.315 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 157.885 36.995 157.955 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 157.605 36.995 157.675 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 173.565 36.995 173.635 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 169.645 36.995 169.715 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 165.725 36.995 165.795 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 161.805 36.995 161.875 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 120.365 36.995 120.435 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 112.525 36.995 112.595 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 108.605 36.995 108.675 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 104.685 36.995 104.755 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 100.765 36.995 100.835 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 96.845 36.995 96.915 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 85.085 36.995 85.155 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 81.165 36.995 81.235 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 77.245 36.995 77.315 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 73.325 36.995 73.395 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 69.405 36.995 69.475 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 65.485 36.995 65.555 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 61.565 36.995 61.635 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 57.645 36.995 57.715 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 53.725 36.995 53.795 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 49.805 36.995 49.875 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 45.885 36.995 45.955 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 41.965 36.995 42.035 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 38.045 36.995 38.115 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 34.125 36.995 34.195 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 30.205 36.995 30.275 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 26.285 36.995 26.355 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 22.365 36.995 22.435 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 18.445 36.995 18.515 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 14.525 36.995 14.595 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 10.605 36.995 10.675 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 6.685 36.995 6.755 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 2.765 36.995 2.835 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 143.885 36.995 143.955 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 152.285 1.715 152.355 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 152.285 2.835 152.355 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.885 0.595 143.955 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.005 0.595 299.075 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 302.925 0.595 302.995 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.045 0.595 143.115 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 302.085 0.595 302.155 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.485 0.595 184.555 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.405 0.595 272.475 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 298.165 0.595 298.235 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 262.885 0.595 262.955 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.365 0.595 239.435 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 215.845 0.595 215.915 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.325 0.595 192.395 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 168.805 0.595 168.875 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 153.405 1.715 153.475 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 153.405 2.835 153.475 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 158.165 37.555 158.235 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.725 0.595 144.795 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p304
    PIN p305
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p306
    PIN p307
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p308
    PIN p309
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p310
    PIN p311
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p312
    PIN p313
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p314
    PIN p315
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p316
    PIN p317
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p318
    PIN p319
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p320
    PIN p321
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p322
    PIN p323
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p324
    PIN p325
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p326
    PIN p327
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p330
    PIN p331
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p332
    PIN p333
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 298.445 0.595 298.515 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.565 0.595 299.635 ;
        END
    END p334
    PIN p335
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 302.365 0.595 302.435 ;
        END
    END p335
    PIN p336
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 155.925 36.995 155.995 ;
        END
    END p336
    PIN p337
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 155.645 0.595 155.715 ;
        END
    END p337
    PIN p338
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 155.085 0.595 155.155 ;
        END
    END p338
    PIN p339
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 153.405 0.595 153.475 ;
        END
    END p339
    PIN p340
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.725 0.595 158.795 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 302.925 36.995 302.995 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 283.325 36.995 283.395 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 279.405 36.995 279.475 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 116.445 36.995 116.515 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 267.645 36.995 267.715 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 263.725 36.995 263.795 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 124.285 36.995 124.355 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 275.485 36.995 275.555 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 271.565 36.995 271.635 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 251.965 36.995 252.035 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 248.045 36.995 248.115 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 259.805 36.995 259.875 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 255.885 36.995 255.955 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 92.925 36.995 92.995 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 89.005 36.995 89.075 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 212.765 36.995 212.835 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 208.845 36.995 208.915 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 220.605 36.995 220.675 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 216.685 36.995 216.755 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 228.445 36.995 228.515 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 224.525 36.995 224.595 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 236.285 36.995 236.355 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 232.365 36.995 232.435 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 244.125 36.995 244.195 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 240.205 36.995 240.275 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 181.405 36.995 181.475 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 177.485 36.995 177.555 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 189.245 36.995 189.315 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 185.325 36.995 185.395 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 197.085 36.995 197.155 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 193.165 36.995 193.235 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 204.925 36.995 204.995 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 201.005 36.995 201.075 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 303.485 0.595 303.555 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 128.205 36.995 128.275 ;
        END
    END p377
    PIN p378
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 132.125 36.995 132.195 ;
        END
    END p378
    PIN p379
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 136.045 36.995 136.115 ;
        END
    END p379
    PIN p380
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 139.965 36.995 140.035 ;
        END
    END p380
    PIN p381
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 287.245 36.995 287.315 ;
        END
    END p381
    PIN p382
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 291.165 36.995 291.235 ;
        END
    END p382
    PIN p383
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 295.085 36.995 295.155 ;
        END
    END p383
    PIN p384
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 299.005 36.995 299.075 ;
        END
    END p384
    PIN p385
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p385
    OBS
      LAYER via2 ;
        RECT  0 0 38.64 307.44 ;
      LAYER metal2 ;
        RECT  0 0 38.64 307.44 ;
      LAYER via1 ;
        RECT  0 0 38.64 307.44 ;
      LAYER metal1 ;
        RECT  0 0 38.64 307.44 ;
    END
END fake_macro_adaptec1_o210920

MACRO fake_macro_adaptec1_o210921
    CLASS BLOCK ;
    SIZE 15.12 BY 275.52 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.725 0.595 137.795 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 140.245 13.475 140.315 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 142.205 13.475 142.275 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 141.925 13.475 141.995 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 57.645 13.475 57.715 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 53.725 13.475 53.795 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 181.405 13.475 181.475 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 146.125 13.475 146.195 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 244.125 13.475 244.195 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 85.085 13.475 85.155 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 208.845 13.475 208.915 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 201.005 13.475 201.075 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 112.525 13.475 112.595 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 22.365 13.475 22.435 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 161.805 13.475 161.875 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 251.965 13.475 252.035 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 255.885 13.475 255.955 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 96.845 13.475 96.915 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 232.365 13.475 232.435 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 259.805 13.475 259.875 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 100.765 13.475 100.835 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 18.445 13.475 18.515 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 77.245 13.475 77.315 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 41.965 13.475 42.035 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 173.565 13.475 173.635 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 157.885 13.475 157.955 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 212.765 13.475 212.835 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 228.445 13.475 228.515 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 89.005 13.475 89.075 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 236.285 13.475 236.355 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 185.325 13.475 185.395 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 104.685 13.475 104.755 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 263.725 13.475 263.795 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 120.365 13.475 120.435 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 193.165 13.475 193.235 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 150.045 13.475 150.115 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.645 13.475 169.715 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 216.685 13.475 216.755 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 189.245 13.475 189.315 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.285 13.475 26.355 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 271.565 13.475 271.635 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 224.525 13.475 224.595 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 248.045 13.475 248.115 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 38.045 13.475 38.115 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 165.725 13.475 165.795 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 240.205 13.475 240.275 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 128.205 13.475 128.275 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 49.805 13.475 49.875 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 197.085 13.475 197.155 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.965 13.475 154.035 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 220.605 13.475 220.675 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 204.925 13.475 204.995 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 177.485 13.475 177.555 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 92.925 13.475 92.995 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 2.765 13.475 2.835 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 6.685 13.475 6.755 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 34.125 13.475 34.195 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 267.645 13.475 267.715 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 45.885 13.475 45.955 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 30.205 13.475 30.275 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 10.605 13.475 10.675 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 65.485 13.475 65.555 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.165 13.475 81.235 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 124.285 13.475 124.355 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 116.445 13.475 116.515 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 61.565 13.475 61.635 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.325 13.475 73.395 ;
        END
    END p68
    PIN p69
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 14.525 13.475 14.595 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 108.605 13.475 108.675 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 69.405 13.475 69.475 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 146.125 0.595 146.195 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 150.045 0.595 150.115 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 153.965 0.595 154.035 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.485 0.595 121.555 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.205 0.595 37.275 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.405 0.595 27.475 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 56.805 0.595 56.875 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 9.765 0.595 9.835 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 146.965 0.595 147.035 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.405 0.595 272.475 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.205 0.595 233.275 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.485 0.595 184.555 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.645 0.595 162.715 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.205 0.595 149.275 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 262.885 0.595 262.955 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 215.845 0.595 215.915 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.325 0.595 192.395 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 168.805 0.595 168.875 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.045 0.595 143.115 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.925 13.475 169.995 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 130.445 13.475 130.515 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 141.645 13.475 141.715 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.605 0.595 136.675 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 145.565 0.595 145.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 146.685 0.595 146.755 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 150.605 0.595 150.675 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 153.405 0.595 153.475 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.525 0.595 154.595 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p303
    PIN p304
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p304
    PIN p305
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p306
    PIN p307
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p308
    PIN p309
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p310
    PIN p311
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p312
    PIN p313
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p314
    PIN p315
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p316
    PIN p317
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p318
    PIN p319
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p320
    PIN p321
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p322
    PIN p323
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p324
    PIN p325
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p326
    PIN p327
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p330
    PIN p331
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p332
    PIN p333
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p334
    PIN p335
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p336
    PIN p337
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p341
    OBS
      LAYER via2 ;
        RECT  0 0 15.12 275.52 ;
      LAYER metal2 ;
        RECT  0 0 15.12 275.52 ;
      LAYER via1 ;
        RECT  0 0 15.12 275.52 ;
      LAYER metal1 ;
        RECT  0 0 15.12 275.52 ;
    END
END fake_macro_adaptec1_o210921

MACRO fake_macro_adaptec1_o210922
    CLASS BLOCK ;
    SIZE 38.64 BY 307.44 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 157.885 36.995 157.955 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 283.325 36.995 283.395 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 279.405 36.995 279.475 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 275.485 36.995 275.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 267.645 36.995 267.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 263.725 36.995 263.795 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 259.805 36.995 259.875 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 255.885 36.995 255.955 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 248.045 36.995 248.115 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 220.605 36.995 220.675 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 197.085 36.995 197.155 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 193.165 36.995 193.235 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 185.325 36.995 185.395 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 181.405 36.995 181.475 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 177.485 36.995 177.555 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 173.565 36.995 173.635 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 169.645 36.995 169.715 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 165.725 36.995 165.795 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 161.805 36.995 161.875 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 104.685 36.995 104.755 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 96.845 36.995 96.915 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 92.925 36.995 92.995 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 85.085 36.995 85.155 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 77.245 36.995 77.315 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 69.405 36.995 69.475 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 65.485 36.995 65.555 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 61.565 36.995 61.635 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 53.725 36.995 53.795 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 41.965 36.995 42.035 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 38.045 36.995 38.115 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 34.125 36.995 34.195 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 30.205 36.995 30.275 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 26.285 36.995 26.355 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 18.445 36.995 18.515 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 14.525 36.995 14.595 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 10.605 36.995 10.675 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 6.685 36.995 6.755 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 2.765 36.995 2.835 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 139.965 36.995 140.035 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 136.045 36.995 136.115 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 132.125 36.995 132.195 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 128.205 36.995 128.275 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 302.925 36.995 302.995 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 143.885 36.995 143.955 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 271.565 36.995 271.635 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 240.205 36.995 240.275 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 236.285 36.995 236.355 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 228.445 36.995 228.515 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 224.525 36.995 224.595 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 216.685 36.995 216.755 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 212.765 36.995 212.835 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 208.845 36.995 208.915 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 204.925 36.995 204.995 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 201.005 36.995 201.075 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 189.245 36.995 189.315 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 124.285 36.995 124.355 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 120.365 36.995 120.435 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 116.445 36.995 116.515 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 112.525 36.995 112.595 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 108.605 36.995 108.675 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 100.765 36.995 100.835 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 89.005 36.995 89.075 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 81.165 36.995 81.235 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 73.325 36.995 73.395 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 57.645 36.995 57.715 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 49.805 36.995 49.875 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 45.885 36.995 45.955 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 22.365 36.995 22.435 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 152.285 1.715 152.355 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 152.285 2.835 152.355 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 152.285 0.595 152.355 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 146.125 36.995 146.195 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 173.845 36.995 173.915 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 147.245 0.595 147.315 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.885 0.595 143.955 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.005 0.595 299.075 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 302.925 0.595 302.995 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.045 0.595 143.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 302.085 0.595 302.155 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.565 0.595 278.635 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.485 0.595 184.555 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.405 0.595 272.475 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 298.165 0.595 298.235 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 262.885 0.595 262.955 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.365 0.595 239.435 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 215.845 0.595 215.915 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.325 0.595 192.395 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 168.805 0.595 168.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 153.405 1.715 153.475 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 153.405 2.835 153.475 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 158.165 37.555 158.235 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.725 0.595 144.795 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p304
    PIN p305
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p306
    PIN p307
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p308
    PIN p309
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p310
    PIN p311
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p312
    PIN p313
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p314
    PIN p315
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p316
    PIN p317
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p318
    PIN p319
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p320
    PIN p321
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p322
    PIN p323
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p324
    PIN p325
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p326
    PIN p327
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p330
    PIN p331
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p332
    PIN p333
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p333
    PIN p334
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p335
    PIN p336
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p337
    PIN p338
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p339
    PIN p340
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p341
    PIN p342
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p343
    PIN p344
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p345
    PIN p346
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p347
    PIN p348
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p349
    PIN p350
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p351
    PIN p352
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p353
    PIN p354
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p355
    PIN p356
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p357
    PIN p358
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p359
    PIN p360
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p361
    PIN p362
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p363
    PIN p364
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p365
    PIN p366
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 298.445 0.595 298.515 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.565 0.595 299.635 ;
        END
    END p367
    PIN p368
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 302.365 0.595 302.435 ;
        END
    END p368
    PIN p369
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 155.925 36.995 155.995 ;
        END
    END p369
    PIN p370
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 155.645 0.595 155.715 ;
        END
    END p370
    PIN p371
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 155.085 0.595 155.155 ;
        END
    END p371
    PIN p372
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 153.405 0.595 153.475 ;
        END
    END p372
    PIN p373
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 157.605 36.995 157.675 ;
        END
    END p373
    PIN p374
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.725 0.595 158.795 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 251.965 36.995 252.035 ;
        END
    END p377
    PIN p378
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 232.365 36.995 232.435 ;
        END
    END p378
    PIN p379
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 244.125 36.995 244.195 ;
        END
    END p379
    PIN p380
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 303.485 0.595 303.555 ;
        END
    END p380
    PIN p381
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 287.245 36.995 287.315 ;
        END
    END p381
    PIN p382
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 291.165 36.995 291.235 ;
        END
    END p382
    PIN p383
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 295.085 36.995 295.155 ;
        END
    END p383
    PIN p384
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 299.005 36.995 299.075 ;
        END
    END p384
    PIN p385
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p385
    OBS
      LAYER via2 ;
        RECT  0 0 38.64 307.44 ;
      LAYER metal2 ;
        RECT  0 0 38.64 307.44 ;
      LAYER via1 ;
        RECT  0 0 38.64 307.44 ;
      LAYER metal1 ;
        RECT  0 0 38.64 307.44 ;
    END
END fake_macro_adaptec1_o210922

MACRO fake_macro_adaptec1_o210923
    CLASS BLOCK ;
    SIZE 15.12 BY 275.52 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 142.205 13.475 142.275 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 57.645 13.475 57.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 53.725 13.475 53.795 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 181.405 13.475 181.475 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 146.125 13.475 146.195 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 244.125 13.475 244.195 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 85.085 13.475 85.155 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 208.845 13.475 208.915 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 201.005 13.475 201.075 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 112.525 13.475 112.595 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 22.365 13.475 22.435 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 161.805 13.475 161.875 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 251.965 13.475 252.035 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 255.885 13.475 255.955 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 96.845 13.475 96.915 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 232.365 13.475 232.435 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 259.805 13.475 259.875 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 100.765 13.475 100.835 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 18.445 13.475 18.515 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 77.245 13.475 77.315 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 41.965 13.475 42.035 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 173.565 13.475 173.635 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 157.885 13.475 157.955 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 212.765 13.475 212.835 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 228.445 13.475 228.515 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 89.005 13.475 89.075 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 236.285 13.475 236.355 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 185.325 13.475 185.395 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 104.685 13.475 104.755 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 263.725 13.475 263.795 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 120.365 13.475 120.435 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 193.165 13.475 193.235 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 150.045 13.475 150.115 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.645 13.475 169.715 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 216.685 13.475 216.755 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 189.245 13.475 189.315 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.285 13.475 26.355 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 271.565 13.475 271.635 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 224.525 13.475 224.595 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 248.045 13.475 248.115 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 38.045 13.475 38.115 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 165.725 13.475 165.795 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 240.205 13.475 240.275 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 128.205 13.475 128.275 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 49.805 13.475 49.875 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 197.085 13.475 197.155 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.965 13.475 154.035 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 220.605 13.475 220.675 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 204.925 13.475 204.995 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 177.485 13.475 177.555 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 92.925 13.475 92.995 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 2.765 13.475 2.835 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 6.685 13.475 6.755 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 34.125 13.475 34.195 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 267.645 13.475 267.715 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 45.885 13.475 45.955 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 30.205 13.475 30.275 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 10.605 13.475 10.675 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 65.485 13.475 65.555 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.165 13.475 81.235 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 124.285 13.475 124.355 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 116.445 13.475 116.515 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 61.565 13.475 61.635 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.325 13.475 73.395 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 14.525 13.475 14.595 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 108.605 13.475 108.675 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 69.405 13.475 69.475 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.725 0.595 137.795 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 140.245 13.475 140.315 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 141.925 13.475 141.995 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 146.125 0.595 146.195 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 150.045 0.595 150.115 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 153.965 0.595 154.035 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.485 0.595 121.555 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.205 0.595 37.275 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.405 0.595 27.475 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.605 0.595 17.675 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 56.805 0.595 56.875 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 9.765 0.595 9.835 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 262.885 0.595 262.955 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 215.845 0.595 215.915 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.325 0.595 192.395 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 168.805 0.595 168.875 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 146.965 0.595 147.035 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.405 0.595 272.475 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.205 0.595 233.275 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.485 0.595 184.555 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.645 0.595 162.715 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.205 0.595 149.275 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.045 0.595 143.115 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.925 13.475 169.995 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 130.445 13.475 130.515 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 141.645 13.475 141.715 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.605 0.595 136.675 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 145.565 0.595 145.635 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 146.685 0.595 146.755 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 150.605 0.595 150.675 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 153.405 0.595 153.475 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.525 0.595 154.595 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p303
    PIN p304
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p304
    PIN p305
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p306
    PIN p307
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p308
    PIN p309
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p310
    PIN p311
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p312
    PIN p313
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p314
    PIN p315
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p316
    PIN p317
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p318
    PIN p319
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p320
    PIN p321
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p322
    PIN p323
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p324
    PIN p325
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p326
    PIN p327
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p330
    PIN p331
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p332
    PIN p333
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p334
    PIN p335
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p336
    PIN p337
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p341
    OBS
      LAYER via2 ;
        RECT  0 0 15.12 275.52 ;
      LAYER metal2 ;
        RECT  0 0 15.12 275.52 ;
      LAYER via1 ;
        RECT  0 0 15.12 275.52 ;
      LAYER metal1 ;
        RECT  0 0 15.12 275.52 ;
    END
END fake_macro_adaptec1_o210923

MACRO fake_macro_adaptec1_o210924
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.685 21.315 181.755 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.405 21.315 153.475 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o210924

MACRO fake_macro_adaptec1_o210925
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.685 21.315 181.755 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.405 21.315 153.475 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p285
    PIN p286
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p287
    PIN p288
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p289
    PIN p290
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p291
    PIN p292
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o210925

MACRO fake_macro_adaptec1_o210926
    CLASS BLOCK ;
    SIZE 38.64 BY 146.16 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 70.245 36.995 70.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 70.525 36.995 70.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 16.205 0.595 16.275 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 20.125 0.595 20.195 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.885 0.595 31.955 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 55.405 0.595 55.475 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 59.325 0.595 59.395 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.125 0.595 83.195 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.045 0.595 87.115 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.885 0.595 94.955 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 98.805 0.595 98.875 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 102.725 0.595 102.795 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.645 0.595 106.715 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.565 0.595 110.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.485 0.595 114.555 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.405 0.595 118.475 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.325 0.595 122.395 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.165 0.595 130.235 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.085 0.595 134.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.005 0.595 138.075 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.925 0.595 141.995 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 97.965 36.995 98.035 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 7.525 36.995 7.595 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 11.445 36.995 11.515 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 15.365 36.995 15.435 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 19.285 36.995 19.355 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 23.205 36.995 23.275 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 27.125 36.995 27.195 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 31.045 36.995 31.115 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 34.965 36.995 35.035 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 38.885 36.995 38.955 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 42.805 36.995 42.875 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 46.725 36.995 46.795 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 50.645 36.995 50.715 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 54.565 36.995 54.635 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 58.485 36.995 58.555 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 62.405 36.995 62.475 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 66.325 36.995 66.395 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 84.245 36.995 84.315 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 88.165 36.995 88.235 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 92.085 36.995 92.155 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 96.005 36.995 96.075 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 99.925 36.995 99.995 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 103.845 36.995 103.915 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 107.765 36.995 107.835 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 111.685 36.995 111.755 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 115.605 36.995 115.675 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 119.525 36.995 119.595 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 123.445 36.995 123.515 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 127.365 36.995 127.435 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 131.285 36.995 131.355 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 135.205 36.995 135.275 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 139.125 36.995 139.195 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 143.045 36.995 143.115 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 3.605 36.995 3.675 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 72.205 36.995 72.275 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.045 0.595 73.115 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.725 0.595 74.795 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 74.725 1.715 74.795 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 74.725 2.835 74.795 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.045 0.595 143.115 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.885 0.595 80.955 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 82.005 36.995 82.075 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  37.485 82.285 37.555 82.355 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 75.845 0.595 75.915 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 75.845 1.715 75.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 75.845 2.835 75.915 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.205 0.595 142.275 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.605 0.595 143.675 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.285 0.595 138.355 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.685 0.595 139.755 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.365 0.595 134.435 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.765 0.595 135.835 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.445 0.595 130.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.845 0.595 131.915 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.525 0.595 126.595 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.925 0.595 127.995 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.605 0.595 122.675 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.005 0.595 124.075 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.685 0.595 118.755 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.085 0.595 120.155 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.765 0.595 114.835 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.845 0.595 110.915 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.245 0.595 112.315 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.925 0.595 106.995 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.325 0.595 108.395 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.005 0.595 103.075 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.405 0.595 104.475 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.085 0.595 99.155 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.485 0.595 100.555 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.165 0.595 95.235 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.565 0.595 96.635 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.245 0.595 91.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.645 0.595 92.715 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.325 0.595 87.395 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.725 0.595 88.795 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.405 0.595 83.475 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.885 0.595 66.955 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.765 0.595 65.835 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.965 0.595 63.035 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.845 0.595 61.915 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 59.045 0.595 59.115 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.925 0.595 57.995 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 55.125 0.595 55.195 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.005 0.595 54.075 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 51.205 0.595 51.275 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.085 0.595 50.155 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.285 0.595 47.355 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.165 0.595 46.235 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.365 0.595 43.435 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.245 0.595 42.315 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.445 0.595 39.515 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.525 0.595 35.595 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.405 0.595 34.475 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.605 0.595 31.675 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.485 0.595 30.555 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.685 0.595 27.755 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.565 0.595 26.635 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.765 0.595 23.835 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.645 0.595 22.715 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.845 0.595 19.915 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.725 0.595 18.795 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.925 0.595 15.995 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.805 0.595 14.875 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 12.005 0.595 12.075 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.885 0.595 10.955 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 8.085 0.595 8.155 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.965 0.595 7.035 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 4.165 0.595 4.235 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.165 0.595 116.235 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.805 0.595 84.875 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.045 0.595 3.115 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.325 0.595 38.395 ;
        END
    END p180
    OBS
      LAYER via2 ;
        RECT  0 0 38.64 146.16 ;
      LAYER metal2 ;
        RECT  0 0 38.64 146.16 ;
      LAYER via1 ;
        RECT  0 0 38.64 146.16 ;
      LAYER metal1 ;
        RECT  0 0 38.64 146.16 ;
    END
END fake_macro_adaptec1_o210926

MACRO fake_macro_adaptec1_o210927
    CLASS BLOCK ;
    SIZE 98 BY 399.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 1.085 90.755 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.885 1.085 87.955 1.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 1.085 86.275 1.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 1.085 84.035 1.155 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 1.085 82.355 1.155 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 1.085 80.675 1.155 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 1.085 78.995 1.155 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 1.085 76.755 1.155 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 1.085 75.075 1.155 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 1.085 68.915 1.155 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 1.085 67.235 1.155 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 1.085 65.555 1.155 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 1.085 63.875 1.155 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 1.085 61.635 1.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.885 1.085 59.955 1.155 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 1.085 58.275 1.155 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 1.085 56.595 1.155 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 1.085 53.235 1.155 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.085 51.555 1.155 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 1.085 49.875 1.155 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 1.085 48.195 1.155 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 1.085 45.955 1.155 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 1.085 44.275 1.155 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 1.085 42.595 1.155 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.845 1.085 40.915 1.155 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 1.085 34.755 1.155 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 1.085 33.075 1.155 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 1.085 30.835 1.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 1.085 29.155 1.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 1.085 27.475 1.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 1.085 25.795 1.155 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 1.085 23.555 1.155 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 1.085 21.875 1.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 21.525 2.835 21.595 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 23.765 3.395 23.835 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 23.765 2.835 23.835 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 26.005 3.395 26.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 28.245 3.395 28.315 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 28.245 2.835 28.315 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 30.485 3.395 30.555 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 30.485 2.835 30.555 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 17.045 3.395 17.115 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 17.045 2.835 17.115 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 19.285 3.395 19.355 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 19.285 2.835 19.355 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.525 3.395 21.595 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 4.725 11.795 4.795 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 4.725 14.595 4.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 4.725 14.035 4.795 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 4.725 15.715 4.795 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.285 1.715 12.355 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 12.285 12.355 12.355 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 11.165 3.395 11.235 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 1.085 91.315 1.155 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 4.725 12.915 4.795 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 11.165 2.835 11.235 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 26.005 2.835 26.075 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 5.845 5.075 5.915 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 5.845 7.315 5.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 1.085 6.195 1.155 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 1.085 11.235 1.155 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 32.445 11.795 32.515 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 49.245 3.395 49.315 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.245 3.395 21.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.765 3.955 30.835 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.205 3.955 30.275 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 28.525 3.955 28.595 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 27.965 3.955 28.035 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 26.285 3.955 26.355 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 25.725 3.955 25.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 24.045 3.955 24.115 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 23.485 3.955 23.555 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 21.805 3.955 21.875 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 1.085 22.435 1.155 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 1.085 24.675 1.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 1.085 26.355 1.155 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 1.085 28.035 1.155 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 1.085 29.715 1.155 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 1.085 31.955 1.155 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 1.085 33.635 1.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 1.085 35.315 1.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 1.085 41.475 1.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 1.085 43.155 1.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 1.085 44.835 1.155 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 1.085 47.075 1.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 1.085 48.755 1.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 1.085 50.435 1.155 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 1.085 52.115 1.155 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 1.085 54.355 1.155 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.085 57.155 1.155 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.085 58.835 1.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 1.085 60.515 1.155 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 1.085 62.755 1.155 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 1.085 64.435 1.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.045 1.085 66.115 1.155 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 1.085 67.795 1.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 1.085 70.035 1.155 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 1.085 75.635 1.155 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 1.085 79.555 1.155 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.165 1.085 81.235 1.155 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 1.085 82.915 1.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 1.085 85.155 1.155 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 1.085 86.835 1.155 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  88.445 1.085 88.515 1.155 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.845 1.715 12.915 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 17.325 91.875 17.395 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 17.325 24.675 17.395 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 17.325 22.995 17.395 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 17.325 47.075 17.395 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 17.325 45.395 17.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 17.325 43.715 17.395 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 17.325 42.035 17.395 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 17.325 35.875 17.395 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 17.325 34.195 17.395 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 17.325 31.955 17.395 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 17.325 30.275 17.395 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 17.325 28.595 17.395 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 17.325 26.915 17.395 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 17.325 66.675 17.395 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 17.325 64.995 17.395 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 17.325 62.755 17.395 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 17.325 61.075 17.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 17.325 59.395 17.395 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 17.325 57.715 17.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 17.325 54.355 17.395 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 17.325 52.675 17.395 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 17.325 50.995 17.395 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 17.325 49.315 17.395 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.565 1.715 12.635 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 19.565 10.115 19.635 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 17.325 89.075 17.395 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 17.325 87.395 17.395 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 17.325 85.155 17.395 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 17.325 83.475 17.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 17.325 81.795 17.395 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 17.325 80.115 17.395 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 17.325 77.875 17.395 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 17.325 76.195 17.395 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 17.325 70.035 17.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 17.325 68.355 17.395 ;
        END
    END p140
    OBS
      LAYER via2 ;
        RECT  0 0 98.14 399.84 ;
      LAYER metal2 ;
        RECT  0 0 98.14 399.84 ;
      LAYER via1 ;
        RECT  0 0 98.14 399.84 ;
      LAYER metal1 ;
        RECT  0 0 98.14 399.84 ;
    END
END fake_macro_adaptec1_o210927

MACRO fake_macro_adaptec1_o210928
    CLASS BLOCK ;
    SIZE 80.08 BY 141.12 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 1.085 76.755 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 1.085 75.075 1.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 1.085 73.395 1.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 1.085 71.715 1.155 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 1.085 69.475 1.155 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 1.085 63.875 1.155 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 1.085 61.635 1.155 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.885 1.085 59.955 1.155 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 1.085 58.275 1.155 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 1.085 56.595 1.155 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 1.085 53.235 1.155 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.085 51.555 1.155 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 1.085 49.875 1.155 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 1.085 48.195 1.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 1.085 45.955 1.155 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 1.085 44.275 1.155 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 1.085 42.595 1.155 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.845 1.085 40.915 1.155 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 1.085 34.755 1.155 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 1.085 33.075 1.155 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 1.085 30.835 1.155 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 1.085 29.155 1.155 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 1.085 27.475 1.155 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 1.085 25.795 1.155 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 1.085 23.555 1.155 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 1.085 21.875 1.155 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 11.165 2.835 11.235 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 26.005 2.835 26.075 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 1.085 6.195 1.155 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 4.725 12.915 4.795 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.525 3.395 21.595 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 19.285 3.395 19.355 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 30.485 3.395 30.555 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 58.205 3.395 58.275 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 28.245 3.395 28.315 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 30.205 3.395 30.275 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 26.005 3.395 26.075 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 27.965 3.395 28.035 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 23.765 3.395 23.835 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 12.285 12.355 12.355 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 11.165 3.395 11.235 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 21.525 2.835 21.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 24.045 3.955 24.115 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 23.765 2.835 23.835 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 26.285 3.955 26.355 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 28.525 3.955 28.595 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 28.245 2.835 28.315 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.765 3.955 30.835 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 30.485 2.835 30.555 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 17.045 3.395 17.115 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 17.045 2.835 17.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 19.565 3.955 19.635 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 19.285 2.835 19.355 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 21.805 3.955 21.875 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 4.725 11.795 4.795 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 4.725 14.595 4.795 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 4.725 14.035 4.795 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 4.725 15.715 4.795 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.285 1.715 12.355 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 5.845 5.075 5.915 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 5.845 7.315 5.915 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 1.085 11.235 1.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 32.445 11.795 32.515 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 1.085 22.435 1.155 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 1.085 24.675 1.155 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 1.085 26.355 1.155 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 1.085 28.035 1.155 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 1.085 29.715 1.155 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 1.085 31.955 1.155 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 1.085 33.635 1.155 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 1.085 35.315 1.155 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 1.085 41.475 1.155 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 1.085 43.155 1.155 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 1.085 44.835 1.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 1.085 47.075 1.155 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 1.085 48.755 1.155 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 1.085 50.435 1.155 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 1.085 52.115 1.155 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 1.085 54.355 1.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.085 57.155 1.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.085 58.835 1.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 1.085 60.515 1.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 1.085 62.755 1.155 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 1.085 64.435 1.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 1.085 70.595 1.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.205 1.085 72.275 1.155 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.885 1.085 73.955 1.155 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 1.085 75.635 1.155 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 17.325 76.195 17.395 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  74.445 17.325 74.515 17.395 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.765 17.325 72.835 17.395 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 17.325 70.595 17.395 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 17.325 64.995 17.395 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 17.325 62.755 17.395 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 17.325 61.075 17.395 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 17.325 59.395 17.395 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 17.325 57.715 17.395 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 17.325 54.355 17.395 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 17.325 30.275 17.395 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 17.325 28.595 17.395 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 17.325 26.915 17.395 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 17.325 24.675 17.395 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 17.325 22.995 17.395 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 17.325 52.675 17.395 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 17.325 50.995 17.395 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 17.325 49.315 17.395 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 17.325 47.075 17.395 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 17.325 45.395 17.395 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 17.325 43.715 17.395 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 17.325 42.035 17.395 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 17.325 35.875 17.395 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 17.325 34.195 17.395 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 17.325 31.955 17.395 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.565 1.715 12.635 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 17.325 77.875 17.395 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.845 1.715 12.915 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 19.565 10.115 19.635 ;
        END
    END p117
    OBS
      LAYER via2 ;
        RECT  0 0 80.08 141.12 ;
      LAYER metal2 ;
        RECT  0 0 80.08 141.12 ;
      LAYER via1 ;
        RECT  0 0 80.08 141.12 ;
      LAYER metal1 ;
        RECT  0 0 80.08 141.12 ;
    END
END fake_macro_adaptec1_o210928

MACRO fake_macro_adaptec1_o210929
    CLASS BLOCK ;
    SIZE 47.6 BY 28.56 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 16.205 1.155 16.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 27.405 14.595 27.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 27.405 10.115 27.475 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 27.405 5.635 27.475 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 26.285 1.155 26.355 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 27.405 15.715 27.475 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 27.405 11.235 27.475 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 27.405 6.755 27.475 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 25.445 1.155 25.515 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.005 1.155 19.075 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 27.405 13.475 27.475 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 27.405 17.955 27.475 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.925 1.155 22.995 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 27.405 7.875 27.475 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 18.725 45.955 18.795 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 10.325 45.955 10.395 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 2.765 22.435 2.835 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.925 27.405 8.995 27.475 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 17.045 45.955 17.115 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 15.365 45.955 15.435 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 13.685 45.955 13.755 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 12.005 45.955 12.075 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 8.645 45.955 8.715 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 6.965 45.955 7.035 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 5.285 45.955 5.355 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 3.605 45.955 3.675 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 27.125 45.955 27.195 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 25.445 45.955 25.515 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 23.765 45.955 23.835 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 22.085 45.955 22.155 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 20.405 45.955 20.475 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 2.765 6.755 2.835 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.085 2.765 15.155 2.835 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 3.045 24.675 3.115 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 2.765 14.035 2.835 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 6.125 13.475 6.195 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 17.885 1.155 17.955 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 14.805 1.155 14.875 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 22.085 1.155 22.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.765 27.405 16.835 27.475 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 27.405 21.875 27.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  20.125 27.405 20.195 27.475 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 2.485 10.115 2.555 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  19.005 2.205 19.075 2.275 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 27.405 12.355 27.475 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  19.005 27.405 19.075 27.475 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 20.125 1.155 20.195 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 27.405 21.315 27.475 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 21.245 1.155 21.315 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 27.405 9.555 27.475 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 27.405 14.035 27.475 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  18.445 27.405 18.515 27.475 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 23.765 1.155 23.835 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 27.405 8.435 27.475 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 27.405 12.915 27.475 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 27.405 17.395 27.475 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 27.405 22.995 27.475 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 2.765 17.395 2.835 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 3.605 11.795 3.675 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 2.765 16.275 2.835 ;
        END
    END p60
    OBS
      LAYER via2 ;
        RECT  0 0 47.6 28.56 ;
      LAYER metal2 ;
        RECT  0 0 47.6 28.56 ;
      LAYER via1 ;
        RECT  0 0 47.6 28.56 ;
      LAYER metal1 ;
        RECT  0 0 47.6 28.56 ;
    END
END fake_macro_adaptec1_o210929

MACRO fake_macro_adaptec1_o210930
    CLASS BLOCK ;
    SIZE 72.24 BY 236.88 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 115.045 68.915 115.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 113.925 69.475 113.995 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.685 0.595 34.755 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 155.925 0.595 155.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.725 0.595 81.795 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.965 0.595 203.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.325 0.595 234.395 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 16.765 0.595 16.835 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 63.805 0.595 63.875 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.845 0.595 110.915 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.325 0.595 136.395 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 152.005 0.595 152.075 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.685 0.595 167.755 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 183.365 0.595 183.435 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 199.045 0.595 199.115 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 214.725 0.595 214.795 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 230.405 0.595 230.475 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 125.405 70.035 125.475 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 153.125 70.035 153.195 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.645 0.595 120.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 119.525 3.955 119.595 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.925 0.595 120.995 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 119.805 70.035 119.875 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 117.845 70.035 117.915 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 115.885 70.035 115.955 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.165 0.595 116.235 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.725 0.595 116.795 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.405 0.595 118.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 117.285 1.155 117.355 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 118.405 3.395 118.475 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 118.405 2.275 118.475 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.645 0.595 218.715 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 187.285 0.595 187.355 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.605 0.595 171.675 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.245 0.595 140.315 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.405 0.595 97.475 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.085 0.595 127.155 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.045 0.595 66.115 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.165 0.595 95.235 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.365 0.595 50.435 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 79.485 0.595 79.555 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.005 0.595 19.075 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.125 0.595 48.195 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.325 0.595 3.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 32.445 0.595 32.515 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.085 0.595 113.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 146.685 0.595 146.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.005 0.595 131.075 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.925 0.595 106.995 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.245 0.595 91.315 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 75.565 0.595 75.635 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 59.885 0.595 59.955 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 44.205 0.595 44.275 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 28.525 0.595 28.595 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 12.845 0.595 12.915 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 113.925 68.355 113.995 ;
        END
    END p77
    PIN p78
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 27.965 70.595 28.035 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 43.645 70.595 43.715 ;
        END
    END p79
    PIN p80
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 59.325 70.595 59.395 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 75.005 70.595 75.075 ;
        END
    END p81
    PIN p82
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 90.685 70.595 90.755 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 106.365 70.595 106.435 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 131.565 70.595 131.635 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 147.245 70.595 147.315 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 162.925 70.595 162.995 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 178.605 70.595 178.675 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 12.285 70.595 12.355 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 194.285 70.595 194.355 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 209.965 70.595 210.035 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 225.645 70.595 225.715 ;
        END
    END p91
    OBS
      LAYER via2 ;
        RECT  0 0 72.24 236.88 ;
      LAYER metal2 ;
        RECT  0 0 72.24 236.88 ;
      LAYER via1 ;
        RECT  0 0 72.24 236.88 ;
      LAYER metal1 ;
        RECT  0 0 72.24 236.88 ;
    END
END fake_macro_adaptec1_o210930

MACRO fake_macro_adaptec1_o210931
    CLASS BLOCK ;
    SIZE 11.2 BY 146.16 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 70.245 9.555 70.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 97.965 9.555 98.035 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.605 0.595 143.675 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 4.165 0.595 4.235 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 16.205 0.595 16.275 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.885 0.595 31.955 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.965 0.595 91.035 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.645 0.595 106.715 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.005 0.595 138.075 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 70.525 9.555 70.595 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 24.045 0.595 24.115 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 51.485 0.595 51.555 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.565 0.595 110.635 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.245 0.595 126.315 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.925 0.595 141.995 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 59.325 0.595 59.395 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.125 0.595 83.195 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.045 0.595 87.115 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 98.805 0.595 98.875 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 102.725 0.595 102.795 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.485 0.595 114.555 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.405 0.595 118.475 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.165 0.595 130.235 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.085 0.595 134.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.045 0.595 143.115 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.685 0.595 139.755 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.205 0.595 142.275 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.765 0.595 135.835 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.285 0.595 138.355 ;
        END
    END p74
    PIN p75
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.845 0.595 131.915 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.365 0.595 134.435 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.925 0.595 127.995 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.445 0.595 130.515 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.005 0.595 124.075 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.525 0.595 126.595 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.085 0.595 120.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.605 0.595 122.675 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.165 0.595 116.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.685 0.595 118.755 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.245 0.595 112.315 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.765 0.595 114.835 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.325 0.595 108.395 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.845 0.595 110.915 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.405 0.595 104.475 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.925 0.595 106.995 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.485 0.595 100.555 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.005 0.595 103.075 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.565 0.595 96.635 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.085 0.595 99.155 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.645 0.595 92.715 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.165 0.595 95.235 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.725 0.595 88.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.245 0.595 91.315 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.805 0.595 84.875 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.325 0.595 87.395 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.765 0.595 65.835 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.405 0.595 83.475 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.845 0.595 61.915 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.885 0.595 66.955 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.925 0.595 57.995 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.965 0.595 63.035 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.005 0.595 54.075 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 59.045 0.595 59.115 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.085 0.595 50.155 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 55.125 0.595 55.195 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.165 0.595 46.235 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 51.205 0.595 51.275 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.245 0.595 42.315 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.285 0.595 47.355 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.325 0.595 38.395 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.365 0.595 43.435 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.405 0.595 34.475 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.445 0.595 39.515 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.485 0.595 30.555 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.525 0.595 35.595 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.565 0.595 26.635 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.605 0.595 31.675 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.645 0.595 22.715 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.685 0.595 27.755 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.725 0.595 18.795 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.765 0.595 23.835 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.805 0.595 14.875 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.845 0.595 19.915 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.885 0.595 10.955 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.925 0.595 15.995 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.965 0.595 7.035 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 12.005 0.595 12.075 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.045 0.595 3.115 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 8.085 0.595 8.155 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 72.205 9.555 72.275 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.045 0.595 73.115 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.885 0.595 80.955 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 82.005 9.555 82.075 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 82.285 10.115 82.355 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 139.125 9.555 139.195 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 143.045 9.555 143.115 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 99.925 9.555 99.995 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 103.845 9.555 103.915 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 107.765 9.555 107.835 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 111.685 9.555 111.755 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 115.605 9.555 115.675 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 119.525 9.555 119.595 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 123.445 9.555 123.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 127.365 9.555 127.435 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 131.285 9.555 131.355 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 135.205 9.555 135.275 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 46.725 9.555 46.795 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 50.645 9.555 50.715 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 54.565 9.555 54.635 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 58.485 9.555 58.555 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 62.405 9.555 62.475 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 66.325 9.555 66.395 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 84.245 9.555 84.315 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 88.165 9.555 88.235 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 92.085 9.555 92.155 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 96.005 9.555 96.075 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 7.525 9.555 7.595 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 11.445 9.555 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 15.365 9.555 15.435 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 19.285 9.555 19.355 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 23.205 9.555 23.275 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 27.125 9.555 27.195 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 31.045 9.555 31.115 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 34.965 9.555 35.035 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 38.885 9.555 38.955 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 42.805 9.555 42.875 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 3.605 9.555 3.675 ;
        END
    END p174
    OBS
      LAYER via2 ;
        RECT  0 0 11.2 146.16 ;
      LAYER metal2 ;
        RECT  0 0 11.2 146.16 ;
      LAYER via1 ;
        RECT  0 0 11.2 146.16 ;
      LAYER metal1 ;
        RECT  0 0 11.2 146.16 ;
    END
END fake_macro_adaptec1_o210931

MACRO fake_macro_adaptec1_o210932
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 51.205 0.595 51.275 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210932

MACRO fake_macro_adaptec1_o210933
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 51.205 0.595 51.275 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210933

MACRO fake_macro_adaptec1_o210934
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 51.205 0.595 51.275 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210934

MACRO fake_macro_adaptec1_o210935
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 51.205 0.595 51.275 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210935

MACRO fake_macro_adaptec1_o210936
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210936

MACRO fake_macro_adaptec1_o210937
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210937

MACRO fake_macro_adaptec1_o210938
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210938

MACRO fake_macro_adaptec1_o210939
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210939

MACRO fake_macro_adaptec1_o210940
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210940

MACRO fake_macro_adaptec1_o210941
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210941

MACRO fake_macro_adaptec1_o210942
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210942

MACRO fake_macro_adaptec1_o210943
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210943

MACRO fake_macro_adaptec1_o210944
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210944

MACRO fake_macro_adaptec1_o210945
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210945

MACRO fake_macro_adaptec1_o210946
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210946

MACRO fake_macro_adaptec1_o210947
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210947

MACRO fake_macro_adaptec1_o210948
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210948

MACRO fake_macro_adaptec1_o210949
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210949

MACRO fake_macro_adaptec1_o210950
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210950

MACRO fake_macro_adaptec1_o210951
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210951

MACRO fake_macro_adaptec1_o210952
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210952

MACRO fake_macro_adaptec1_o210953
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210953

MACRO fake_macro_adaptec1_o210954
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210954

MACRO fake_macro_adaptec1_o210955
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210955

MACRO fake_macro_adaptec1_o210956
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210956

MACRO fake_macro_adaptec1_o210957
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210957

MACRO fake_macro_adaptec1_o210958
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210958

MACRO fake_macro_adaptec1_o210959
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210959

MACRO fake_macro_adaptec1_o210960
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o210960

MACRO fake_macro_adaptec1_o210961
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210961

MACRO fake_macro_adaptec1_o210962
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210962

MACRO fake_macro_adaptec1_o210963
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210963

MACRO fake_macro_adaptec1_o210964
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210964

MACRO fake_macro_adaptec1_o210965
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210965

MACRO fake_macro_adaptec1_o210966
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210966

MACRO fake_macro_adaptec1_o210967
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210967

MACRO fake_macro_adaptec1_o210968
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210968

MACRO fake_macro_adaptec1_o210969
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210969

MACRO fake_macro_adaptec1_o210970
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210970

MACRO fake_macro_adaptec1_o210971
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210971

MACRO fake_macro_adaptec1_o210972
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210972

MACRO fake_macro_adaptec1_o210973
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210973

MACRO fake_macro_adaptec1_o210974
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210974

MACRO fake_macro_adaptec1_o210975
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210975

MACRO fake_macro_adaptec1_o210976
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210976

MACRO fake_macro_adaptec1_o210977
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210977

MACRO fake_macro_adaptec1_o210978
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210978

MACRO fake_macro_adaptec1_o210979
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210979

MACRO fake_macro_adaptec1_o210980
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210980

MACRO fake_macro_adaptec1_o210981
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210981

MACRO fake_macro_adaptec1_o210982
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210982

MACRO fake_macro_adaptec1_o210983
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210983

MACRO fake_macro_adaptec1_o210984
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210984

MACRO fake_macro_adaptec1_o210985
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210985

MACRO fake_macro_adaptec1_o210986
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210986

MACRO fake_macro_adaptec1_o210987
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210987

MACRO fake_macro_adaptec1_o210988
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210988

MACRO fake_macro_adaptec1_o210989
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210989

MACRO fake_macro_adaptec1_o210990
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210990

MACRO fake_macro_adaptec1_o210991
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210991

MACRO fake_macro_adaptec1_o210992
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210992

MACRO fake_macro_adaptec1_o210993
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210993

MACRO fake_macro_adaptec1_o210994
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210994

MACRO fake_macro_adaptec1_o210995
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210995

MACRO fake_macro_adaptec1_o210996
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210996

MACRO fake_macro_adaptec1_o210997
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210997

MACRO fake_macro_adaptec1_o210998
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210998

MACRO fake_macro_adaptec1_o210999
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o210999

MACRO fake_macro_adaptec1_o211000
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211000

MACRO fake_macro_adaptec1_o211001
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211001

MACRO fake_macro_adaptec1_o211002
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211002

MACRO fake_macro_adaptec1_o211003
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211003

MACRO fake_macro_adaptec1_o211004
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211004

MACRO fake_macro_adaptec1_o211005
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211005

MACRO fake_macro_adaptec1_o211006
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211006

MACRO fake_macro_adaptec1_o211007
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211007

MACRO fake_macro_adaptec1_o211008
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211008

MACRO fake_macro_adaptec1_o211009
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211009

MACRO fake_macro_adaptec1_o211010
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211010

MACRO fake_macro_adaptec1_o211011
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211011

MACRO fake_macro_adaptec1_o211012
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211012

MACRO fake_macro_adaptec1_o211013
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211013

MACRO fake_macro_adaptec1_o211014
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211014

MACRO fake_macro_adaptec1_o211015
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211015

MACRO fake_macro_adaptec1_o211016
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211016

MACRO fake_macro_adaptec1_o211017
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211017

MACRO fake_macro_adaptec1_o211018
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211018

MACRO fake_macro_adaptec1_o211019
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211019

MACRO fake_macro_adaptec1_o211020
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211020

MACRO fake_macro_adaptec1_o211021
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211021

MACRO fake_macro_adaptec1_o211022
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211022

MACRO fake_macro_adaptec1_o211023
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211023

MACRO fake_macro_adaptec1_o211024
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211024

MACRO fake_macro_adaptec1_o211025
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211025

MACRO fake_macro_adaptec1_o211026
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211026

MACRO fake_macro_adaptec1_o211027
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211027

MACRO fake_macro_adaptec1_o211028
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211028

MACRO fake_macro_adaptec1_o211029
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211029

MACRO fake_macro_adaptec1_o211030
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211030

MACRO fake_macro_adaptec1_o211031
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211031

MACRO fake_macro_adaptec1_o211032
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211032

MACRO fake_macro_adaptec1_o211033
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211033

MACRO fake_macro_adaptec1_o211034
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211034

MACRO fake_macro_adaptec1_o211035
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211035

MACRO fake_macro_adaptec1_o211036
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211036

MACRO fake_macro_adaptec1_o211037
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211037

MACRO fake_macro_adaptec1_o211038
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211038

MACRO fake_macro_adaptec1_o211039
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211039

MACRO fake_macro_adaptec1_o211040
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211040

MACRO fake_macro_adaptec1_o211041
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211041

MACRO fake_macro_adaptec1_o211042
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211042

MACRO fake_macro_adaptec1_o211043
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211043

MACRO fake_macro_adaptec1_o211044
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211044

MACRO fake_macro_adaptec1_o211045
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211045

MACRO fake_macro_adaptec1_o211046
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 3.325 58.835 3.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 7.805 58.835 7.875 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 8.085 58.835 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.365 58.275 8.435 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 3.885 56.595 3.955 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211046

MACRO fake_macro_adaptec1_o211047
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211047

MACRO fake_macro_adaptec1_o211048
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211048

MACRO fake_macro_adaptec1_o211049
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211049

MACRO fake_macro_adaptec1_o211050
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 3.325 58.835 3.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 8.085 58.835 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 7.805 58.835 7.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.365 58.275 8.435 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 3.885 56.595 3.955 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211050

MACRO fake_macro_adaptec1_o211051
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211051

MACRO fake_macro_adaptec1_o211052
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211052

MACRO fake_macro_adaptec1_o211053
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 8.085 58.835 8.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 3.325 58.835 3.395 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 7.805 58.835 7.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.365 58.275 8.435 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 3.885 56.595 3.955 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211053

MACRO fake_macro_adaptec1_o211054
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211054

MACRO fake_macro_adaptec1_o211055
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 3.325 58.835 3.395 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 8.085 58.835 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 7.805 58.835 7.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.365 58.275 8.435 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 3.885 56.595 3.955 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211055

MACRO fake_macro_adaptec1_o211056
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 8.085 58.835 8.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 3.325 58.835 3.395 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 7.805 58.835 7.875 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.365 58.275 8.435 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 3.885 56.595 3.955 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211056

MACRO fake_macro_adaptec1_o211057
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211057

MACRO fake_macro_adaptec1_o211058
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211058

MACRO fake_macro_adaptec1_o211059
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211059

MACRO fake_macro_adaptec1_o211060
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211060

MACRO fake_macro_adaptec1_o211061
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211061

MACRO fake_macro_adaptec1_o211062
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211062

MACRO fake_macro_adaptec1_o211063
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211063

MACRO fake_macro_adaptec1_o211064
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211064

MACRO fake_macro_adaptec1_o211065
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211065

MACRO fake_macro_adaptec1_o211066
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211066

MACRO fake_macro_adaptec1_o211067
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211067

MACRO fake_macro_adaptec1_o211068
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211068

MACRO fake_macro_adaptec1_o211069
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211069

MACRO fake_macro_adaptec1_o211070
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211070

MACRO fake_macro_adaptec1_o211071
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211071

MACRO fake_macro_adaptec1_o211072
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211072

MACRO fake_macro_adaptec1_o211073
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211073

MACRO fake_macro_adaptec1_o211074
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211074

MACRO fake_macro_adaptec1_o211075
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211075

MACRO fake_macro_adaptec1_o211076
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211076

MACRO fake_macro_adaptec1_o211077
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211077

MACRO fake_macro_adaptec1_o211078
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211078

MACRO fake_macro_adaptec1_o211079
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211079

MACRO fake_macro_adaptec1_o211080
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211080

MACRO fake_macro_adaptec1_o211081
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211081

MACRO fake_macro_adaptec1_o211082
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211082

MACRO fake_macro_adaptec1_o211083
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211083

MACRO fake_macro_adaptec1_o211084
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211084

MACRO fake_macro_adaptec1_o211085
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211085

MACRO fake_macro_adaptec1_o211086
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211086

MACRO fake_macro_adaptec1_o211087
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211087

MACRO fake_macro_adaptec1_o211088
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211088

MACRO fake_macro_adaptec1_o211089
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211089

MACRO fake_macro_adaptec1_o211090
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211090

MACRO fake_macro_adaptec1_o211091
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211091

MACRO fake_macro_adaptec1_o211092
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211092

MACRO fake_macro_adaptec1_o211093
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211093

MACRO fake_macro_adaptec1_o211094
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211094

MACRO fake_macro_adaptec1_o211095
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211095

MACRO fake_macro_adaptec1_o211096
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211096

MACRO fake_macro_adaptec1_o211097
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211097

MACRO fake_macro_adaptec1_o211098
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211098

MACRO fake_macro_adaptec1_o211099
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211099

MACRO fake_macro_adaptec1_o211100
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211100

MACRO fake_macro_adaptec1_o211101
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211101

MACRO fake_macro_adaptec1_o211102
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211102

MACRO fake_macro_adaptec1_o211103
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211103

MACRO fake_macro_adaptec1_o211104
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211104

MACRO fake_macro_adaptec1_o211105
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211105

MACRO fake_macro_adaptec1_o211106
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211106

MACRO fake_macro_adaptec1_o211107
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211107

MACRO fake_macro_adaptec1_o211108
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211108

MACRO fake_macro_adaptec1_o211109
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211109

MACRO fake_macro_adaptec1_o211110
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211110

MACRO fake_macro_adaptec1_o211111
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211111

MACRO fake_macro_adaptec1_o211112
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211112

MACRO fake_macro_adaptec1_o211113
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211113

MACRO fake_macro_adaptec1_o211114
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211114

MACRO fake_macro_adaptec1_o211115
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211115

MACRO fake_macro_adaptec1_o211116
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211116

MACRO fake_macro_adaptec1_o211117
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211117

MACRO fake_macro_adaptec1_o211118
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211118

MACRO fake_macro_adaptec1_o211119
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211119

MACRO fake_macro_adaptec1_o211120
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211120

MACRO fake_macro_adaptec1_o211121
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211121

MACRO fake_macro_adaptec1_o211122
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211122

MACRO fake_macro_adaptec1_o211123
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211123

MACRO fake_macro_adaptec1_o211124
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.645 1.155 1.715 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.925 1.155 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 5.845 3.395 5.915 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211124

MACRO fake_macro_adaptec1_o211125
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211125

MACRO fake_macro_adaptec1_o211126
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211126

MACRO fake_macro_adaptec1_o211127
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211127

MACRO fake_macro_adaptec1_o211128
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.645 1.155 1.715 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.925 1.155 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 5.845 3.395 5.915 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211128

MACRO fake_macro_adaptec1_o211129
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211129

MACRO fake_macro_adaptec1_o211130
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211130

MACRO fake_macro_adaptec1_o211131
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211131

MACRO fake_macro_adaptec1_o211132
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211132

MACRO fake_macro_adaptec1_o211133
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211133

MACRO fake_macro_adaptec1_o211134
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211134

MACRO fake_macro_adaptec1_o211135
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211135

MACRO fake_macro_adaptec1_o211136
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211136

MACRO fake_macro_adaptec1_o211137
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211137

MACRO fake_macro_adaptec1_o211138
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211138

MACRO fake_macro_adaptec1_o211139
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211139

MACRO fake_macro_adaptec1_o211140
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211140

MACRO fake_macro_adaptec1_o211141
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211141

MACRO fake_macro_adaptec1_o211142
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211142

MACRO fake_macro_adaptec1_o211143
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211143

MACRO fake_macro_adaptec1_o211144
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211144

MACRO fake_macro_adaptec1_o211145
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211145

MACRO fake_macro_adaptec1_o211146
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211146

MACRO fake_macro_adaptec1_o211147
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211147

MACRO fake_macro_adaptec1_o211148
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211148

MACRO fake_macro_adaptec1_o211149
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211149

MACRO fake_macro_adaptec1_o211150
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211150

MACRO fake_macro_adaptec1_o211151
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211151

MACRO fake_macro_adaptec1_o211152
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211152

MACRO fake_macro_adaptec1_o211153
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.645 1.155 1.715 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.925 1.155 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 5.845 3.395 5.915 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211153

MACRO fake_macro_adaptec1_o211154
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211154

MACRO fake_macro_adaptec1_o211155
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211155

MACRO fake_macro_adaptec1_o211156
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211156

MACRO fake_macro_adaptec1_o211157
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211157

MACRO fake_macro_adaptec1_o211158
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211158

MACRO fake_macro_adaptec1_o211159
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211159

MACRO fake_macro_adaptec1_o211160
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211160

MACRO fake_macro_adaptec1_o211161
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211161

MACRO fake_macro_adaptec1_o211162
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211162

MACRO fake_macro_adaptec1_o211163
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211163

MACRO fake_macro_adaptec1_o211164
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211164

MACRO fake_macro_adaptec1_o211165
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211165

MACRO fake_macro_adaptec1_o211166
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211166

MACRO fake_macro_adaptec1_o211167
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211167

MACRO fake_macro_adaptec1_o211168
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211168

MACRO fake_macro_adaptec1_o211169
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211169

MACRO fake_macro_adaptec1_o211170
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211170

MACRO fake_macro_adaptec1_o211171
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211171

MACRO fake_macro_adaptec1_o211172
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211172

MACRO fake_macro_adaptec1_o211173
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211173

MACRO fake_macro_adaptec1_o211174
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211174

MACRO fake_macro_adaptec1_o211175
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211175

MACRO fake_macro_adaptec1_o211176
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211176

MACRO fake_macro_adaptec1_o211177
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211177

MACRO fake_macro_adaptec1_o211178
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211178

MACRO fake_macro_adaptec1_o211179
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211179

MACRO fake_macro_adaptec1_o211180
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211180

MACRO fake_macro_adaptec1_o211181
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211181

MACRO fake_macro_adaptec1_o211182
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211182

MACRO fake_macro_adaptec1_o211183
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211183

MACRO fake_macro_adaptec1_o211184
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211184

MACRO fake_macro_adaptec1_o211185
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211185

MACRO fake_macro_adaptec1_o211186
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211186

MACRO fake_macro_adaptec1_o211187
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211187

MACRO fake_macro_adaptec1_o211188
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211188

MACRO fake_macro_adaptec1_o211189
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211189

MACRO fake_macro_adaptec1_o211190
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211190

MACRO fake_macro_adaptec1_o211191
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211191

MACRO fake_macro_adaptec1_o211192
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211192

MACRO fake_macro_adaptec1_o211193
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211193

MACRO fake_macro_adaptec1_o211194
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211194

MACRO fake_macro_adaptec1_o211195
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211195

MACRO fake_macro_adaptec1_o211196
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 3.325 5.075 3.395 ;
        END
    END p2
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211196

MACRO fake_macro_adaptec1_o211197
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.365 57.155 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 5.285 56.595 5.355 ;
        END
    END p2
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211197

MACRO fake_macro_adaptec1_o211198
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 58.765 5.635 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211198

MACRO fake_macro_adaptec1_o211199
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 58.765 5.635 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211199

MACRO fake_macro_adaptec1_o211200
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 6.685 57.155 6.755 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 3.325 58.275 3.395 ;
        END
    END p3
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211200

MACRO fake_macro_adaptec1_o211201
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211201

MACRO fake_macro_adaptec1_o211202
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211202

MACRO fake_macro_adaptec1_o211203
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211203

MACRO fake_macro_adaptec1_o211204
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211204

MACRO fake_macro_adaptec1_o211205
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211205

MACRO fake_macro_adaptec1_o211206
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211206

MACRO fake_macro_adaptec1_o211207
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211207

MACRO fake_macro_adaptec1_o211208
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211208

MACRO fake_macro_adaptec1_o211209
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211209

MACRO fake_macro_adaptec1_o211210
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211210

MACRO fake_macro_adaptec1_o211211
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211211

MACRO fake_macro_adaptec1_o211212
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211212

MACRO fake_macro_adaptec1_o211213
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211213

MACRO fake_macro_adaptec1_o211214
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211214

MACRO fake_macro_adaptec1_o211215
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211215

MACRO fake_macro_adaptec1_o211216
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211216

MACRO fake_macro_adaptec1_o211217
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211217

MACRO fake_macro_adaptec1_o211218
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211218

MACRO fake_macro_adaptec1_o211219
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211219

MACRO fake_macro_adaptec1_o211220
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211220

MACRO fake_macro_adaptec1_o211221
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211221

MACRO fake_macro_adaptec1_o211222
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211222

MACRO fake_macro_adaptec1_o211223
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211223

MACRO fake_macro_adaptec1_o211224
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211224

MACRO fake_macro_adaptec1_o211225
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211225

MACRO fake_macro_adaptec1_o211226
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211226

MACRO fake_macro_adaptec1_o211227
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211227

MACRO fake_macro_adaptec1_o211228
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211228

MACRO fake_macro_adaptec1_o211229
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211229

MACRO fake_macro_adaptec1_o211230
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211230

MACRO fake_macro_adaptec1_o211231
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211231

MACRO fake_macro_adaptec1_o211232
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211232

MACRO fake_macro_adaptec1_o211233
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211233

MACRO fake_macro_adaptec1_o211234
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211234

MACRO fake_macro_adaptec1_o211235
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211235

MACRO fake_macro_adaptec1_o211236
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211236

MACRO fake_macro_adaptec1_o211237
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211237

MACRO fake_macro_adaptec1_o211238
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211238

MACRO fake_macro_adaptec1_o211239
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211239

MACRO fake_macro_adaptec1_o211240
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211240

MACRO fake_macro_adaptec1_o211241
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211241

MACRO fake_macro_adaptec1_o211242
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211242

MACRO fake_macro_adaptec1_o211243
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211243

MACRO fake_macro_adaptec1_o211244
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211244

MACRO fake_macro_adaptec1_o211245
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211245

MACRO fake_macro_adaptec1_o211246
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211246

MACRO fake_macro_adaptec1_o211247
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211247

MACRO fake_macro_adaptec1_o211248
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211248

MACRO fake_macro_adaptec1_o211249
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211249

MACRO fake_macro_adaptec1_o211250
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211250

MACRO fake_macro_adaptec1_o211251
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211251

MACRO fake_macro_adaptec1_o211252
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211252

MACRO fake_macro_adaptec1_o211253
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211253

MACRO fake_macro_adaptec1_o211254
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211254

MACRO fake_macro_adaptec1_o211255
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211255

MACRO fake_macro_adaptec1_o211256
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211256

MACRO fake_macro_adaptec1_o211257
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211257

MACRO fake_macro_adaptec1_o211258
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211258

MACRO fake_macro_adaptec1_o211259
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211259

MACRO fake_macro_adaptec1_o211260
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211260

MACRO fake_macro_adaptec1_o211261
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211261

MACRO fake_macro_adaptec1_o211262
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211262

MACRO fake_macro_adaptec1_o211263
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211263

MACRO fake_macro_adaptec1_o211264
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211264

MACRO fake_macro_adaptec1_o211265
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211265

MACRO fake_macro_adaptec1_o211266
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211266

MACRO fake_macro_adaptec1_o211267
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211267

MACRO fake_macro_adaptec1_o211268
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211268

MACRO fake_macro_adaptec1_o211269
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211269

MACRO fake_macro_adaptec1_o211270
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211270

MACRO fake_macro_adaptec1_o211271
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211271

MACRO fake_macro_adaptec1_o211272
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211272

MACRO fake_macro_adaptec1_o211273
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211273

MACRO fake_macro_adaptec1_o211274
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211274

MACRO fake_macro_adaptec1_o211275
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211275

MACRO fake_macro_adaptec1_o211276
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211276

MACRO fake_macro_adaptec1_o211277
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211277

MACRO fake_macro_adaptec1_o211278
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211278

MACRO fake_macro_adaptec1_o211279
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211279

MACRO fake_macro_adaptec1_o211280
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211280

MACRO fake_macro_adaptec1_o211281
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211281

MACRO fake_macro_adaptec1_o211282
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211282

MACRO fake_macro_adaptec1_o211283
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211283

MACRO fake_macro_adaptec1_o211284
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211284

MACRO fake_macro_adaptec1_o211285
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211285

MACRO fake_macro_adaptec1_o211286
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211286

MACRO fake_macro_adaptec1_o211287
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211287

MACRO fake_macro_adaptec1_o211288
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211288

MACRO fake_macro_adaptec1_o211289
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211289

MACRO fake_macro_adaptec1_o211290
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211290

MACRO fake_macro_adaptec1_o211291
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211291

MACRO fake_macro_adaptec1_o211292
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211292

MACRO fake_macro_adaptec1_o211293
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211293

MACRO fake_macro_adaptec1_o211294
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211294

MACRO fake_macro_adaptec1_o211295
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211295

MACRO fake_macro_adaptec1_o211296
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211296

MACRO fake_macro_adaptec1_o211297
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211297

MACRO fake_macro_adaptec1_o211298
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211298

MACRO fake_macro_adaptec1_o211299
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211299

MACRO fake_macro_adaptec1_o211300
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211300

MACRO fake_macro_adaptec1_o211301
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211301

MACRO fake_macro_adaptec1_o211302
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211302

MACRO fake_macro_adaptec1_o211303
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211303

MACRO fake_macro_adaptec1_o211304
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211304

MACRO fake_macro_adaptec1_o211305
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211305

MACRO fake_macro_adaptec1_o211306
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211306

MACRO fake_macro_adaptec1_o211307
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211307

MACRO fake_macro_adaptec1_o211308
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211308

MACRO fake_macro_adaptec1_o211309
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211309

MACRO fake_macro_adaptec1_o211310
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211310

MACRO fake_macro_adaptec1_o211311
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211311

MACRO fake_macro_adaptec1_o211312
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211312

MACRO fake_macro_adaptec1_o211313
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211313

MACRO fake_macro_adaptec1_o211314
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211314

MACRO fake_macro_adaptec1_o211315
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211315

MACRO fake_macro_adaptec1_o211316
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211316

MACRO fake_macro_adaptec1_o211317
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211317

MACRO fake_macro_adaptec1_o211318
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211318

MACRO fake_macro_adaptec1_o211319
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211319

MACRO fake_macro_adaptec1_o211320
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211320

MACRO fake_macro_adaptec1_o211321
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211321

MACRO fake_macro_adaptec1_o211322
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211322

MACRO fake_macro_adaptec1_o211323
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211323

MACRO fake_macro_adaptec1_o211324
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211324

MACRO fake_macro_adaptec1_o211325
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211325

MACRO fake_macro_adaptec1_o211326
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211326

MACRO fake_macro_adaptec1_o211327
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211327

MACRO fake_macro_adaptec1_o211328
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211328

MACRO fake_macro_adaptec1_o211329
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211329

MACRO fake_macro_adaptec1_o211330
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211330

MACRO fake_macro_adaptec1_o211331
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211331

MACRO fake_macro_adaptec1_o211332
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211332

MACRO fake_macro_adaptec1_o211333
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211333

MACRO fake_macro_adaptec1_o211334
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211334

MACRO fake_macro_adaptec1_o211335
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211335

MACRO fake_macro_adaptec1_o211336
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211336

MACRO fake_macro_adaptec1_o211337
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211337

MACRO fake_macro_adaptec1_o211338
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211338

MACRO fake_macro_adaptec1_o211339
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211339

MACRO fake_macro_adaptec1_o211340
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211340

MACRO fake_macro_adaptec1_o211341
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211341

MACRO fake_macro_adaptec1_o211342
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211342

MACRO fake_macro_adaptec1_o211343
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211343

MACRO fake_macro_adaptec1_o211344
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.645 1.155 1.715 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.925 1.155 1.995 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 5.845 3.395 5.915 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211344

MACRO fake_macro_adaptec1_o211345
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211345

MACRO fake_macro_adaptec1_o211346
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211346

MACRO fake_macro_adaptec1_o211347
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211347

MACRO fake_macro_adaptec1_o211348
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.645 1.155 1.715 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 6.405 1.155 6.475 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 1.925 1.155 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 5.845 3.395 5.915 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211348

MACRO fake_macro_adaptec1_o211349
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211349

MACRO fake_macro_adaptec1_o211350
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211350

MACRO fake_macro_adaptec1_o211351
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211351

MACRO fake_macro_adaptec1_o211352
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211352

MACRO fake_macro_adaptec1_o211353
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211353

MACRO fake_macro_adaptec1_o211354
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211354

MACRO fake_macro_adaptec1_o211355
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211355

MACRO fake_macro_adaptec1_o211356
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211356

MACRO fake_macro_adaptec1_o211357
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211357

MACRO fake_macro_adaptec1_o211358
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211358

MACRO fake_macro_adaptec1_o211359
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p5
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211359

MACRO fake_macro_adaptec1_o211360
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211360

MACRO fake_macro_adaptec1_o211361
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211361

MACRO fake_macro_adaptec1_o211362
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211362

MACRO fake_macro_adaptec1_o211363
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211363

MACRO fake_macro_adaptec1_o211364
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p1
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211364

MACRO fake_macro_adaptec1_o211365
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211365

MACRO fake_macro_adaptec1_o211366
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211366

MACRO fake_macro_adaptec1_o211367
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211367

MACRO fake_macro_adaptec1_o211368
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211368

MACRO fake_macro_adaptec1_o211369
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211369

MACRO fake_macro_adaptec1_o211370
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211370

MACRO fake_macro_adaptec1_o211371
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211371

MACRO fake_macro_adaptec1_o211372
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211372

MACRO fake_macro_adaptec1_o211373
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p3
    PIN p4
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p4
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211373

MACRO fake_macro_adaptec1_o211374
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.765 1.715 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 58.765 6.195 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 60.165 1.715 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.205 1.155 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.565 56.805 5.635 56.875 ;
        END
    END p6
    PIN p7
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p7
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211374

MACRO fake_macro_adaptec1_o211375
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211375

MACRO fake_macro_adaptec1_o211376
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211376

MACRO fake_macro_adaptec1_o211377
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211377

MACRO fake_macro_adaptec1_o211378
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211378

MACRO fake_macro_adaptec1_o211379
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211379

MACRO fake_macro_adaptec1_o211380
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211380

MACRO fake_macro_adaptec1_o211381
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211381

MACRO fake_macro_adaptec1_o211382
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211382

MACRO fake_macro_adaptec1_o211383
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211383

MACRO fake_macro_adaptec1_o211384
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211384

MACRO fake_macro_adaptec1_o211385
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211385

MACRO fake_macro_adaptec1_o211386
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211386

MACRO fake_macro_adaptec1_o211387
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211387

MACRO fake_macro_adaptec1_o211388
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211388

MACRO fake_macro_adaptec1_o211389
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211389

MACRO fake_macro_adaptec1_o211390
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211390

MACRO fake_macro_adaptec1_o211391
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211391

MACRO fake_macro_adaptec1_o211392
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211392

MACRO fake_macro_adaptec1_o211393
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211393

MACRO fake_macro_adaptec1_o211394
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211394

MACRO fake_macro_adaptec1_o211395
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211395

MACRO fake_macro_adaptec1_o211396
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 58.765 2.835 58.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 58.765 7.315 58.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 58.765 7.875 58.835 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 60.165 2.835 60.235 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 58.205 1.715 58.275 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 56.805 1.155 56.875 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  -0.035 18.165 0.035 18.235 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211396

MACRO fake_macro_adaptec1_o211397
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211397

MACRO fake_macro_adaptec1_o211398
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211398

MACRO fake_macro_adaptec1_o211399
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211399

MACRO fake_macro_adaptec1_o211400
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211400

MACRO fake_macro_adaptec1_o211401
    CLASS BLOCK ;
    SIZE 10.08 BY 60.48 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 1.365 6.755 1.435 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.365 2.275 1.435 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.365 1.715 1.435 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.685 29.085 6.755 29.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.805 1.925 7.875 1.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  8.365 3.325 8.435 3.395 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal2 ;
        RECT  0 0 10.08 60.48 ;
      LAYER via1 ;
        RECT  0 0 10.08 60.48 ;
      LAYER metal1 ;
        RECT  0 0 10.08 60.48 ;
    END
END fake_macro_adaptec1_o211401

MACRO fake_macro_adaptec1_o211402
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211402

MACRO fake_macro_adaptec1_o211403
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 2.765 1.155 2.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 7.525 1.155 7.595 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 8.085 1.155 8.155 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 1.645 1.715 1.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.045 1.155 3.115 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 1.365 3.395 1.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 -0.035 42.035 0.035 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211403

MACRO fake_macro_adaptec1_o211404
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211404

MACRO fake_macro_adaptec1_o211405
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211405

MACRO fake_macro_adaptec1_o211406
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211406

MACRO fake_macro_adaptec1_o211407
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211407

MACRO fake_macro_adaptec1_o211408
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211408

MACRO fake_macro_adaptec1_o211409
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211409

MACRO fake_macro_adaptec1_o211410
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211410

MACRO fake_macro_adaptec1_o211411
    CLASS BLOCK ;
    SIZE 60.48 BY 10.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.965 58.835 7.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 2.205 58.835 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.645 58.835 1.715 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 6.685 58.835 6.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 8.085 58.275 8.155 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 8.365 56.595 8.435 ;
        END
    END p5
    PIN p6
        DIRECTION INOUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 9.765 17.955 9.835 ;
        END
    END p6
    OBS
      LAYER via2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal2 ;
        RECT  0 0 60.48 10.08 ;
      LAYER via1 ;
        RECT  0 0 60.48 10.08 ;
      LAYER metal1 ;
        RECT  0 0 60.48 10.08 ;
    END
END fake_macro_adaptec1_o211411

MACRO fake_macro_adaptec1_o211412
    CLASS BLOCK ;
    SIZE 110.88 BY 141.12 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 139.685 11.235 139.755 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 129.605 2.835 129.675 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 119.245 2.835 119.315 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 117.005 3.395 117.075 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 117.005 2.835 117.075 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 114.765 3.395 114.835 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 114.765 2.835 114.835 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 112.525 3.395 112.595 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 112.525 2.835 112.595 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 110.285 3.395 110.355 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 110.285 2.835 110.355 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 123.725 3.395 123.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 123.725 2.835 123.795 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 121.485 3.395 121.555 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 121.485 2.835 121.555 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 119.245 3.395 119.315 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 136.045 11.795 136.115 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 136.045 14.595 136.115 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 136.045 14.035 136.115 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 136.045 15.715 136.115 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 128.485 1.715 128.555 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 134.925 7.315 134.995 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 139.685 6.195 139.755 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 140.805 11.795 140.875 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 128.205 1.715 128.275 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 121.205 10.115 121.275 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 136.045 12.915 136.115 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 127.925 1.715 127.995 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 139.685 21.875 139.755 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 139.685 23.555 139.755 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 139.685 25.795 139.755 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 139.685 27.475 139.755 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 139.685 29.155 139.755 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 139.685 30.835 139.755 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 139.685 33.075 139.755 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 139.685 34.755 139.755 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.845 139.685 40.915 139.755 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 139.685 42.595 139.755 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 139.685 44.275 139.755 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 139.685 45.955 139.755 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 139.685 48.195 139.755 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 139.685 49.875 139.755 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 139.685 51.555 139.755 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 139.685 53.235 139.755 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 139.685 56.595 139.755 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 139.685 58.275 139.755 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.885 139.685 59.955 139.755 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 139.685 61.635 139.755 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 139.685 63.875 139.755 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 139.685 65.555 139.755 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 139.685 67.235 139.755 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 139.685 68.915 139.755 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 139.685 75.075 139.755 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 139.685 76.755 139.755 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 139.685 78.995 139.755 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 139.685 80.675 139.755 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 139.685 82.355 139.755 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 139.685 84.035 139.755 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 139.685 86.275 139.755 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.885 139.685 87.955 139.755 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 139.685 90.755 139.755 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  92.365 139.685 92.435 139.755 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 139.685 94.675 139.755 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 139.685 96.355 139.755 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 139.685 102.515 139.755 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.125 139.685 104.195 139.755 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  105.805 139.685 105.875 139.755 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  107.485 139.685 107.555 139.755 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 134.925 5.075 134.995 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 139.685 22.435 139.755 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 139.685 24.675 139.755 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 139.685 26.355 139.755 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 139.685 28.035 139.755 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 139.685 29.715 139.755 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 139.685 31.955 139.755 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 139.685 33.635 139.755 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 139.685 35.315 139.755 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 139.685 41.475 139.755 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 139.685 43.155 139.755 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 139.685 44.835 139.755 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 139.685 47.075 139.755 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 139.685 48.755 139.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 139.685 50.435 139.755 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 139.685 52.115 139.755 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 139.685 54.355 139.755 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 139.685 57.155 139.755 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 139.685 58.835 139.755 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 139.685 60.515 139.755 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 139.685 62.755 139.755 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 139.685 64.435 139.755 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.045 139.685 66.115 139.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 139.685 67.795 139.755 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.685 70.035 139.755 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 139.685 75.635 139.755 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 139.685 77.875 139.755 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 139.685 79.555 139.755 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.165 139.685 81.235 139.755 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 139.685 82.915 139.755 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 139.685 85.155 139.755 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 139.685 86.835 139.755 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  88.445 139.685 88.515 139.755 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 139.685 91.315 139.755 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 139.685 93.555 139.755 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 139.685 95.235 139.755 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 139.685 96.915 139.755 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 139.685 103.075 139.755 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.685 139.685 104.755 139.755 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.365 139.685 106.435 139.755 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  108.605 139.685 108.675 139.755 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 128.485 12.355 128.555 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 140.805 3.395 140.875 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 121.765 3.955 121.835 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 110.565 3.955 110.635 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 110.005 3.955 110.075 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 112.805 3.955 112.875 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 112.245 3.955 112.315 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 115.045 3.955 115.115 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 114.485 3.955 114.555 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 117.285 3.955 117.355 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 129.605 3.395 129.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 123.445 43.715 123.515 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 123.445 42.035 123.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 123.445 35.875 123.515 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 123.445 34.195 123.515 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 123.445 31.955 123.515 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 123.445 30.275 123.515 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 123.445 28.595 123.515 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 123.445 26.915 123.515 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 123.445 24.675 123.515 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 123.445 22.995 123.515 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 123.445 62.755 123.515 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 123.445 61.075 123.515 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 123.445 59.395 123.515 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 123.445 57.715 123.515 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 123.445 54.355 123.515 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 123.445 52.675 123.515 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 123.445 50.995 123.515 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 123.445 49.315 123.515 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 123.445 47.075 123.515 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 123.445 45.395 123.515 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 123.445 85.155 123.515 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 123.445 83.475 123.515 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 123.445 81.795 123.515 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 123.445 80.115 123.515 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 123.445 77.875 123.515 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 123.445 76.195 123.515 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 123.445 70.035 123.515 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 123.445 68.355 123.515 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 123.445 66.675 123.515 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 123.445 64.995 123.515 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  108.605 123.445 108.675 123.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.925 123.445 106.995 123.515 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  105.245 123.445 105.315 123.515 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.565 123.445 103.635 123.515 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 123.445 97.475 123.515 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 123.445 95.795 123.515 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 123.445 93.555 123.515 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 123.445 91.875 123.515 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 123.445 89.075 123.515 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 123.445 87.395 123.515 ;
        END
    END p159
    OBS
      LAYER via2 ;
        RECT  0 0 110.88 141.12 ;
      LAYER metal2 ;
        RECT  0 0 110.88 141.12 ;
      LAYER via1 ;
        RECT  0 0 110.88 141.12 ;
      LAYER metal1 ;
        RECT  0 0 110.88 141.12 ;
    END
END fake_macro_adaptec1_o211412

MACRO fake_macro_adaptec1_o211413
    CLASS BLOCK ;
    SIZE 110.88 BY 141.12 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.165 1.085 11.235 1.155 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 11.165 2.835 11.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 21.525 2.835 21.595 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 23.765 3.395 23.835 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 23.765 2.835 23.835 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 26.005 3.395 26.075 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 26.005 2.835 26.075 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 28.245 3.395 28.315 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 28.245 2.835 28.315 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 30.485 3.395 30.555 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 30.485 2.835 30.555 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 17.045 3.395 17.115 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 17.045 2.835 17.115 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 19.285 3.395 19.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 19.285 2.835 19.355 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.525 3.395 21.595 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 4.725 11.795 4.795 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  14.525 4.725 14.595 4.795 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 4.725 14.035 4.795 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  15.645 4.725 15.715 4.795 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.285 1.715 12.355 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  7.245 5.845 7.315 5.915 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  6.125 1.085 6.195 1.155 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 32.445 11.795 32.515 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.565 1.715 12.635 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 19.565 10.115 19.635 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.845 4.725 12.915 4.795 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 12.845 1.715 12.915 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  5.005 5.845 5.075 5.915 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 1.085 21.875 1.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  23.485 1.085 23.555 1.155 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  25.725 1.085 25.795 1.155 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.405 1.085 27.475 1.155 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.085 1.085 29.155 1.155 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.765 1.085 30.835 1.155 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.005 1.085 33.075 1.155 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.685 1.085 34.755 1.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  40.845 1.085 40.915 1.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  42.525 1.085 42.595 1.155 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.205 1.085 44.275 1.155 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.885 1.085 45.955 1.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.125 1.085 48.195 1.155 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.805 1.085 49.875 1.155 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  51.485 1.085 51.555 1.155 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  53.165 1.085 53.235 1.155 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  56.525 1.085 56.595 1.155 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.205 1.085 58.275 1.155 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.885 1.085 59.955 1.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.565 1.085 61.635 1.155 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 1.085 63.875 1.155 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 1.085 65.555 1.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 1.085 67.235 1.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 1.085 68.915 1.155 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 1.085 75.075 1.155 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 1.085 76.755 1.155 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 1.085 78.995 1.155 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 1.085 80.675 1.155 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 1.085 82.355 1.155 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.965 1.085 84.035 1.155 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.205 1.085 86.275 1.155 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.885 1.085 87.955 1.155 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  90.685 1.085 90.755 1.155 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  92.365 1.085 92.435 1.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  94.605 1.085 94.675 1.155 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 1.085 96.355 1.155 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  102.445 1.085 102.515 1.155 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.125 1.085 104.195 1.155 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  105.805 1.085 105.875 1.155 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  107.485 1.085 107.555 1.155 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.365 1.085 22.435 1.155 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 1.085 24.675 1.155 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.285 1.085 26.355 1.155 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  27.965 1.085 28.035 1.155 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  29.645 1.085 29.715 1.155 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 1.085 31.955 1.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  33.565 1.085 33.635 1.155 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.245 1.085 35.315 1.155 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.405 1.085 41.475 1.155 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.085 1.085 43.155 1.155 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  44.765 1.085 44.835 1.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 1.085 47.075 1.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  48.685 1.085 48.755 1.155 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.365 1.085 50.435 1.155 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.045 1.085 52.115 1.155 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 1.085 54.355 1.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.085 1.085 57.155 1.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  58.765 1.085 58.835 1.155 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  60.445 1.085 60.515 1.155 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 1.085 62.755 1.155 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 1.085 64.435 1.155 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.045 1.085 66.115 1.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 1.085 67.795 1.155 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 1.085 70.035 1.155 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 1.085 75.635 1.155 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 1.085 77.875 1.155 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 1.085 79.555 1.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.165 1.085 81.235 1.155 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.845 1.085 82.915 1.155 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 1.085 85.155 1.155 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  86.765 1.085 86.835 1.155 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  88.445 1.085 88.515 1.155 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.245 1.085 91.315 1.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 1.085 93.555 1.155 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.165 1.085 95.235 1.155 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 1.085 96.915 1.155 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.005 1.085 103.075 1.155 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  104.685 1.085 104.755 1.155 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.365 1.085 106.435 1.155 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  108.605 1.085 108.675 1.155 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  12.285 12.285 12.355 12.355 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 49.245 3.395 49.315 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 21.245 3.395 21.315 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.765 3.955 30.835 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 30.205 3.955 30.275 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 28.525 3.955 28.595 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 27.965 3.955 28.035 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 26.285 3.955 26.355 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 25.725 3.955 25.795 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 24.045 3.955 24.115 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 11.165 3.395 11.235 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  47.005 17.325 47.075 17.395 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  45.325 17.325 45.395 17.395 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  85.085 17.325 85.155 17.395 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  83.405 17.325 83.475 17.395 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 17.325 81.795 17.395 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 17.325 80.115 17.395 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 17.325 77.875 17.395 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 17.325 76.195 17.395 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 17.325 70.035 17.395 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 17.325 68.355 17.395 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 17.325 66.675 17.395 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 17.325 64.995 17.395 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  108.605 17.325 108.675 17.395 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  106.925 17.325 106.995 17.395 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  105.245 17.325 105.315 17.395 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  103.565 17.325 103.635 17.395 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 17.325 97.475 17.395 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  95.725 17.325 95.795 17.395 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  93.485 17.325 93.555 17.395 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  91.805 17.325 91.875 17.395 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  89.005 17.325 89.075 17.395 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  87.325 17.325 87.395 17.395 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  43.645 17.325 43.715 17.395 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  41.965 17.325 42.035 17.395 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  35.805 17.325 35.875 17.395 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  34.125 17.325 34.195 17.395 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  31.885 17.325 31.955 17.395 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  30.205 17.325 30.275 17.395 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  28.525 17.325 28.595 17.395 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  26.845 17.325 26.915 17.395 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  24.605 17.325 24.675 17.395 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  22.925 17.325 22.995 17.395 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  62.685 17.325 62.755 17.395 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  61.005 17.325 61.075 17.395 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  59.325 17.325 59.395 17.395 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  57.645 17.325 57.715 17.395 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  54.285 17.325 54.355 17.395 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  52.605 17.325 52.675 17.395 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  50.925 17.325 50.995 17.395 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  49.245 17.325 49.315 17.395 ;
        END
    END p159
    OBS
      LAYER via2 ;
        RECT  0 0 110.88 141.12 ;
      LAYER metal2 ;
        RECT  0 0 110.88 141.12 ;
      LAYER via1 ;
        RECT  0 0 110.88 141.12 ;
      LAYER metal1 ;
        RECT  0 0 110.88 141.12 ;
    END
END fake_macro_adaptec1_o211413

MACRO fake_macro_adaptec1_o211414
    CLASS BLOCK ;
    SIZE 19.6 BY 304.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 158.165 17.395 158.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 300.685 0.595 300.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 157.045 17.395 157.115 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 156.765 0.595 156.835 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 156.205 0.595 156.275 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 159.845 0.595 159.915 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.405 0.595 160.475 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 142.205 17.395 142.275 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 169.925 17.395 169.995 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 145.005 0.595 145.075 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.845 0.595 271.915 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.765 0.595 275.835 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 285.285 0.595 285.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 281.365 0.595 281.435 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.845 0.595 173.915 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.685 0.595 167.755 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.165 0.595 137.235 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.925 0.595 267.995 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 265.685 0.595 265.755 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 246.085 0.595 246.155 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.325 0.595 234.395 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.885 0.595 220.955 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 199.045 0.595 199.115 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.605 0.595 185.675 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.085 0.595 162.155 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.445 0.595 291.515 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.245 0.595 252.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 238.245 0.595 238.315 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.205 0.595 205.275 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.605 0.595 171.675 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.725 0.595 228.795 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.805 0.595 224.875 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.645 0.595 218.715 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.045 0.595 213.115 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.125 0.595 209.195 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.285 0.595 201.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.445 0.595 193.515 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 191.205 0.595 191.275 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.685 0.595 181.755 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 179.445 0.595 179.515 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.085 0.595 260.155 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.165 0.595 256.235 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.325 0.595 248.395 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.485 0.595 240.555 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.285 0.595 299.355 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.365 0.595 295.435 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.525 0.595 287.595 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 163.485 0.595 163.555 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.405 0.595 167.475 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.325 0.595 171.395 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 175.245 0.595 175.315 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 179.165 0.595 179.235 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 183.085 0.595 183.155 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 187.005 0.595 187.075 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.925 0.595 190.995 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.845 0.595 194.915 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 198.765 0.595 198.835 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.685 0.595 202.755 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 206.605 0.595 206.675 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 210.525 0.595 210.595 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 214.445 0.595 214.515 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.365 0.595 218.435 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 222.285 0.595 222.355 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 226.205 0.595 226.275 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 230.125 0.595 230.195 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.045 0.595 234.115 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 237.965 0.595 238.035 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.885 0.595 241.955 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 245.805 0.595 245.875 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 249.725 0.595 249.795 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 253.645 0.595 253.715 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 257.565 0.595 257.635 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 261.485 0.595 261.555 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 265.405 0.595 265.475 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 269.325 0.595 269.395 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 273.245 0.595 273.315 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 277.165 0.595 277.235 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 281.085 0.595 281.155 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 285.005 0.595 285.075 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.925 0.595 288.995 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.845 0.595 292.915 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 296.765 0.595 296.835 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.565 0.595 299.635 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 152.285 17.395 152.355 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.445 0.595 151.515 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 150.885 0.595 150.955 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 152.285 0.595 152.355 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 159.005 16.275 159.075 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 186.725 16.275 186.795 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.925 0.595 162.995 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.765 0.595 170.835 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.685 0.595 174.755 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.605 0.595 178.675 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.525 0.595 182.595 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.445 0.595 186.515 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.365 0.595 190.435 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 198.205 0.595 198.275 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.125 0.595 202.195 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.965 0.595 210.035 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.885 0.595 213.955 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.805 0.595 217.875 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.725 0.595 221.795 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.645 0.595 225.715 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.565 0.595 229.635 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.485 0.595 233.555 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 237.405 0.595 237.475 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.325 0.595 241.395 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 245.245 0.595 245.315 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 249.165 0.595 249.235 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 253.085 0.595 253.155 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 257.005 0.595 257.075 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.925 0.595 260.995 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.845 0.595 264.915 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.765 0.595 268.835 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.845 0.595 166.915 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.285 0.595 194.355 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 206.045 0.595 206.115 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.365 0.595 288.435 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.685 0.595 272.755 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.285 0.595 292.355 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.605 0.595 276.675 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 296.205 0.595 296.275 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.525 0.595 280.595 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 300.125 0.595 300.195 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.445 0.595 284.515 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 265.405 17.955 265.475 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 85.085 17.395 85.155 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 81.165 17.395 81.235 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 77.245 17.395 77.315 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 73.325 17.395 73.395 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 69.405 17.395 69.475 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 65.485 17.395 65.555 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 61.565 17.395 61.635 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 57.645 17.395 57.715 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 53.725 17.395 53.795 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 49.805 17.395 49.875 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 45.885 17.395 45.955 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 41.965 17.395 42.035 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 38.045 17.395 38.115 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 34.125 17.395 34.195 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 30.205 17.395 30.275 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 26.285 17.395 26.355 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 22.365 17.395 22.435 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 18.445 17.395 18.515 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 14.525 17.395 14.595 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 10.605 17.395 10.675 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 6.685 17.395 6.755 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 2.765 17.395 2.835 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 300.125 17.395 300.195 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 296.205 17.395 296.275 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 292.285 17.395 292.355 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 288.365 17.395 288.435 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 284.445 17.395 284.515 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 280.525 17.395 280.595 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 276.605 17.395 276.675 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 272.685 17.395 272.755 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 268.765 17.395 268.835 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 264.845 17.395 264.915 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 45.325 17.955 45.395 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 41.405 17.955 41.475 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 37.485 17.955 37.555 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 33.565 17.955 33.635 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 29.645 17.955 29.715 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 25.725 17.955 25.795 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 21.805 17.955 21.875 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 17.885 17.955 17.955 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 13.965 17.955 14.035 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 10.045 17.955 10.115 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 260.925 17.395 260.995 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 257.005 17.395 257.075 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 253.085 17.395 253.155 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 249.165 17.395 249.235 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 245.245 17.395 245.315 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 241.325 17.395 241.395 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 237.405 17.395 237.475 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 84.525 17.955 84.595 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 233.485 17.395 233.555 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 80.605 17.955 80.675 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 229.565 17.395 229.635 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 76.685 17.955 76.755 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 225.645 17.395 225.715 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 72.765 17.955 72.835 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 68.845 17.955 68.915 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 64.925 17.955 64.995 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 61.005 17.955 61.075 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 57.085 17.955 57.155 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 53.165 17.955 53.235 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 49.245 17.955 49.315 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 221.725 17.395 221.795 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 217.805 17.395 217.875 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 213.885 17.395 213.955 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 209.965 17.395 210.035 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 206.045 17.395 206.115 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 202.125 17.395 202.195 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 198.205 17.395 198.275 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 194.285 17.395 194.355 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 190.365 17.395 190.435 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 186.445 17.395 186.515 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 182.525 17.395 182.595 ;
        END
    END p377
    PIN p378
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 178.605 17.395 178.675 ;
        END
    END p378
    PIN p379
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 174.685 17.395 174.755 ;
        END
    END p379
    PIN p380
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 170.765 17.395 170.835 ;
        END
    END p380
    PIN p381
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 166.845 17.395 166.915 ;
        END
    END p381
    PIN p382
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 162.925 17.395 162.995 ;
        END
    END p382
    PIN p383
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 139.965 17.395 140.035 ;
        END
    END p383
    PIN p384
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 6.125 17.955 6.195 ;
        END
    END p384
    PIN p385
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 136.045 17.395 136.115 ;
        END
    END p385
    PIN p386
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 2.205 17.955 2.275 ;
        END
    END p386
    PIN p387
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 132.125 17.395 132.195 ;
        END
    END p387
    PIN p388
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 128.205 17.395 128.275 ;
        END
    END p388
    PIN p389
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 124.285 17.395 124.355 ;
        END
    END p389
    PIN p390
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 120.365 17.395 120.435 ;
        END
    END p390
    PIN p391
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 116.445 17.395 116.515 ;
        END
    END p391
    PIN p392
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 112.525 17.395 112.595 ;
        END
    END p392
    PIN p393
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 108.605 17.395 108.675 ;
        END
    END p393
    PIN p394
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 104.685 17.395 104.755 ;
        END
    END p394
    PIN p395
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 100.765 17.395 100.835 ;
        END
    END p395
    PIN p396
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 222.285 17.955 222.355 ;
        END
    END p396
    PIN p397
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 96.845 17.395 96.915 ;
        END
    END p397
    PIN p398
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 218.365 17.955 218.435 ;
        END
    END p398
    PIN p399
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 92.925 17.395 92.995 ;
        END
    END p399
    PIN p400
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 214.445 17.955 214.515 ;
        END
    END p400
    PIN p401
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 89.005 17.395 89.075 ;
        END
    END p401
    PIN p402
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 210.525 17.955 210.595 ;
        END
    END p402
    PIN p403
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 206.605 17.955 206.675 ;
        END
    END p403
    PIN p404
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 202.685 17.955 202.755 ;
        END
    END p404
    PIN p405
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 198.765 17.955 198.835 ;
        END
    END p405
    PIN p406
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 194.845 17.955 194.915 ;
        END
    END p406
    PIN p407
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 190.925 17.955 190.995 ;
        END
    END p407
    PIN p408
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 187.005 17.955 187.075 ;
        END
    END p408
    PIN p409
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 261.485 17.955 261.555 ;
        END
    END p409
    PIN p410
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 257.565 17.955 257.635 ;
        END
    END p410
    PIN p411
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 253.645 17.955 253.715 ;
        END
    END p411
    PIN p412
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 249.725 17.955 249.795 ;
        END
    END p412
    PIN p413
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 245.805 17.955 245.875 ;
        END
    END p413
    PIN p414
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 241.885 17.955 241.955 ;
        END
    END p414
    PIN p415
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 237.965 17.955 238.035 ;
        END
    END p415
    PIN p416
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 234.045 17.955 234.115 ;
        END
    END p416
    PIN p417
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 230.125 17.955 230.195 ;
        END
    END p417
    PIN p418
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 226.205 17.955 226.275 ;
        END
    END p418
    PIN p419
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 123.725 17.955 123.795 ;
        END
    END p419
    PIN p420
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 119.805 17.955 119.875 ;
        END
    END p420
    PIN p421
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 115.885 17.955 115.955 ;
        END
    END p421
    PIN p422
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 111.965 17.955 112.035 ;
        END
    END p422
    PIN p423
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 108.045 17.955 108.115 ;
        END
    END p423
    PIN p424
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 104.125 17.955 104.195 ;
        END
    END p424
    PIN p425
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 100.205 17.955 100.275 ;
        END
    END p425
    PIN p426
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 96.285 17.955 96.355 ;
        END
    END p426
    PIN p427
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 92.365 17.955 92.435 ;
        END
    END p427
    PIN p428
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 88.445 17.955 88.515 ;
        END
    END p428
    PIN p429
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 183.085 17.955 183.155 ;
        END
    END p429
    PIN p430
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 179.165 17.955 179.235 ;
        END
    END p430
    PIN p431
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 175.245 17.955 175.315 ;
        END
    END p431
    PIN p432
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 171.325 17.955 171.395 ;
        END
    END p432
    PIN p433
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 167.405 17.955 167.475 ;
        END
    END p433
    PIN p434
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 163.485 17.955 163.555 ;
        END
    END p434
    PIN p435
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 139.405 17.955 139.475 ;
        END
    END p435
    PIN p436
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 135.485 17.955 135.555 ;
        END
    END p436
    PIN p437
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 131.565 17.955 131.635 ;
        END
    END p437
    PIN p438
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 300.685 17.955 300.755 ;
        END
    END p438
    PIN p439
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 127.645 17.955 127.715 ;
        END
    END p439
    PIN p440
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 296.765 17.955 296.835 ;
        END
    END p440
    PIN p441
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 292.845 17.955 292.915 ;
        END
    END p441
    PIN p442
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 288.925 17.955 288.995 ;
        END
    END p442
    PIN p443
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 285.005 17.955 285.075 ;
        END
    END p443
    PIN p444
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 281.085 17.955 281.155 ;
        END
    END p444
    PIN p445
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 277.165 17.955 277.235 ;
        END
    END p445
    PIN p446
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 273.245 17.955 273.315 ;
        END
    END p446
    PIN p447
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 269.325 17.955 269.395 ;
        END
    END p447
    OBS
      LAYER via2 ;
        RECT  0 0 19.6 304.08 ;
      LAYER metal2 ;
        RECT  0 0 19.6 304.08 ;
      LAYER via1 ;
        RECT  0 0 19.6 304.08 ;
      LAYER metal1 ;
        RECT  0 0 19.6 304.08 ;
    END
END fake_macro_adaptec1_o211414

MACRO fake_macro_adaptec1_o211415
    CLASS BLOCK ;
    SIZE 15.12 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.805 0.595 252.875 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.205 0.595 233.275 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.325 0.595 178.395 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.725 0.595 158.795 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.085 0.595 141.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.485 0.595 121.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.965 13.475 154.035 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.685 13.475 153.755 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 152.005 13.475 152.075 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 181.685 13.475 181.755 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 142.205 13.475 142.275 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.405 13.475 153.475 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 295.085 13.475 295.155 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 291.165 13.475 291.235 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 287.245 13.475 287.315 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 283.325 13.475 283.395 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 279.405 13.475 279.475 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 275.485 13.475 275.555 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 271.565 13.475 271.635 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 267.645 13.475 267.715 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 263.725 13.475 263.795 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 259.805 13.475 259.875 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 85.085 13.475 85.155 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.165 13.475 81.235 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 77.245 13.475 77.315 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.325 13.475 73.395 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 69.405 13.475 69.475 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 65.485 13.475 65.555 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 61.565 13.475 61.635 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 57.645 13.475 57.715 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 53.725 13.475 53.795 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 49.805 13.475 49.875 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 45.885 13.475 45.955 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 41.965 13.475 42.035 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 38.045 13.475 38.115 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 34.125 13.475 34.195 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 30.205 13.475 30.275 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.285 13.475 26.355 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 22.365 13.475 22.435 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 18.445 13.475 18.515 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 14.525 13.475 14.595 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 10.605 13.475 10.675 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 6.685 13.475 6.755 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 2.765 13.475 2.835 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 255.885 13.475 255.955 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 251.965 13.475 252.035 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 248.045 13.475 248.115 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 244.125 13.475 244.195 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 240.205 13.475 240.275 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 236.285 13.475 236.355 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 232.365 13.475 232.435 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 228.445 13.475 228.515 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 224.525 13.475 224.595 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 220.605 13.475 220.675 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 216.685 13.475 216.755 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 212.765 13.475 212.835 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 208.845 13.475 208.915 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 204.925 13.475 204.995 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 201.005 13.475 201.075 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 197.085 13.475 197.155 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 193.165 13.475 193.235 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 189.245 13.475 189.315 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 185.325 13.475 185.395 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 181.405 13.475 181.475 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 177.485 13.475 177.555 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 173.565 13.475 173.635 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.645 13.475 169.715 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 165.725 13.475 165.795 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 161.805 13.475 161.875 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 157.885 13.475 157.955 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 139.965 13.475 140.035 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 136.045 13.475 136.115 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 132.125 13.475 132.195 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 128.205 13.475 128.275 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 124.285 13.475 124.355 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 120.365 13.475 120.435 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 116.445 13.475 116.515 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 112.525 13.475 112.595 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 108.605 13.475 108.675 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 104.685 13.475 104.755 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 100.765 13.475 100.835 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 96.845 13.475 96.915 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 92.925 13.475 92.995 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 89.005 13.475 89.075 ;
        END
    END p371
    OBS
      LAYER via2 ;
        RECT  0 0 15.12 299.04 ;
      LAYER metal2 ;
        RECT  0 0 15.12 299.04 ;
      LAYER via1 ;
        RECT  0 0 15.12 299.04 ;
      LAYER metal1 ;
        RECT  0 0 15.12 299.04 ;
    END
END fake_macro_adaptec1_o211415

MACRO fake_macro_adaptec1_o211416
    CLASS BLOCK ;
    SIZE 19.6 BY 304.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 158.165 17.395 158.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 300.685 0.595 300.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 157.045 17.395 157.115 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 156.765 0.595 156.835 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 156.205 0.595 156.275 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 159.845 0.595 159.915 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 142.205 17.395 142.275 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 169.925 17.395 169.995 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 145.005 0.595 145.075 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.765 0.595 275.835 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 281.365 0.595 281.435 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.845 0.595 271.915 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.325 0.595 248.395 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.885 0.595 220.955 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 199.045 0.595 199.115 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 179.445 0.595 179.515 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.525 0.595 287.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.165 0.595 256.235 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.725 0.595 228.795 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.205 0.595 205.275 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.605 0.595 185.675 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.085 0.595 162.155 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.165 0.595 137.235 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.805 0.595 224.875 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.645 0.595 218.715 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.045 0.595 213.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.125 0.595 209.195 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.285 0.595 201.355 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.445 0.595 193.515 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 191.205 0.595 191.275 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.685 0.595 181.755 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.845 0.595 173.915 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.605 0.595 171.675 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.685 0.595 167.755 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.925 0.595 267.995 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 265.685 0.595 265.755 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.085 0.595 260.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.245 0.595 252.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 246.085 0.595 246.155 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.485 0.595 240.555 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 238.245 0.595 238.315 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.325 0.595 234.395 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.285 0.595 299.355 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.365 0.595 295.435 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.445 0.595 291.515 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 152.285 17.395 152.355 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.445 0.595 151.515 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 150.885 0.595 150.955 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 152.285 0.595 152.355 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 159.005 16.275 159.075 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.925 0.595 162.995 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.765 0.595 170.835 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.685 0.595 174.755 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.605 0.595 178.675 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.525 0.595 182.595 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.445 0.595 186.515 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.365 0.595 190.435 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 198.205 0.595 198.275 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.125 0.595 202.195 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.965 0.595 210.035 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.885 0.595 213.955 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.805 0.595 217.875 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.725 0.595 221.795 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.645 0.595 225.715 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.565 0.595 229.635 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.485 0.595 233.555 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 237.405 0.595 237.475 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.325 0.595 241.395 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 245.245 0.595 245.315 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 249.165 0.595 249.235 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 253.085 0.595 253.155 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 257.005 0.595 257.075 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.925 0.595 260.995 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.845 0.595 264.915 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.765 0.595 268.835 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.845 0.595 166.915 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.285 0.595 194.355 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 206.045 0.595 206.115 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.365 0.595 288.435 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.685 0.595 272.755 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.285 0.595 292.355 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.605 0.595 276.675 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 296.205 0.595 296.275 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.525 0.595 280.595 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 300.125 0.595 300.195 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.445 0.595 284.515 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.405 0.595 160.475 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 285.285 0.595 285.355 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 163.485 0.595 163.555 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.405 0.595 167.475 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.325 0.595 171.395 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 175.245 0.595 175.315 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 179.165 0.595 179.235 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 183.085 0.595 183.155 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 187.005 0.595 187.075 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.925 0.595 190.995 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.845 0.595 194.915 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 198.765 0.595 198.835 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.685 0.595 202.755 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 206.605 0.595 206.675 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 210.525 0.595 210.595 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 214.445 0.595 214.515 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.365 0.595 218.435 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 222.285 0.595 222.355 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 226.205 0.595 226.275 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 230.125 0.595 230.195 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.045 0.595 234.115 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 237.965 0.595 238.035 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.885 0.595 241.955 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 245.805 0.595 245.875 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 249.725 0.595 249.795 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 253.645 0.595 253.715 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 257.565 0.595 257.635 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 261.485 0.595 261.555 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 265.405 0.595 265.475 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 269.325 0.595 269.395 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 273.245 0.595 273.315 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 277.165 0.595 277.235 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 281.085 0.595 281.155 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 285.005 0.595 285.075 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.925 0.595 288.995 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.845 0.595 292.915 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 296.765 0.595 296.835 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.565 0.595 299.635 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 186.725 16.275 186.795 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 85.085 17.395 85.155 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 81.165 17.395 81.235 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 77.245 17.395 77.315 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 73.325 17.395 73.395 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 69.405 17.395 69.475 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 65.485 17.395 65.555 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 61.565 17.395 61.635 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 57.645 17.395 57.715 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 53.725 17.395 53.795 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 49.805 17.395 49.875 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 45.885 17.395 45.955 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 41.965 17.395 42.035 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 38.045 17.395 38.115 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 34.125 17.395 34.195 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 30.205 17.395 30.275 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 26.285 17.395 26.355 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 22.365 17.395 22.435 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 18.445 17.395 18.515 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 14.525 17.395 14.595 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 10.605 17.395 10.675 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 6.685 17.395 6.755 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 2.765 17.395 2.835 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 45.325 17.955 45.395 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 41.405 17.955 41.475 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 37.485 17.955 37.555 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 33.565 17.955 33.635 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 29.645 17.955 29.715 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 300.125 17.395 300.195 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 25.725 17.955 25.795 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 296.205 17.395 296.275 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 21.805 17.955 21.875 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 292.285 17.395 292.355 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 17.885 17.955 17.955 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 260.925 17.395 260.995 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 288.365 17.395 288.435 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 13.965 17.955 14.035 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 257.005 17.395 257.075 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 284.445 17.395 284.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 10.045 17.955 10.115 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 253.085 17.395 253.155 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 280.525 17.395 280.595 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 249.165 17.395 249.235 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 276.605 17.395 276.675 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 245.245 17.395 245.315 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 272.685 17.395 272.755 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 241.325 17.395 241.395 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 268.765 17.395 268.835 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 237.405 17.395 237.475 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 264.845 17.395 264.915 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 233.485 17.395 233.555 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 229.565 17.395 229.635 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 84.525 17.955 84.595 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 225.645 17.395 225.715 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 80.605 17.955 80.675 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 76.685 17.955 76.755 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 72.765 17.955 72.835 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 68.845 17.955 68.915 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 64.925 17.955 64.995 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 61.005 17.955 61.075 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 57.085 17.955 57.155 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 221.725 17.395 221.795 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 53.165 17.955 53.235 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 217.805 17.395 217.875 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 49.245 17.955 49.315 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 213.885 17.395 213.955 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 209.965 17.395 210.035 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 206.045 17.395 206.115 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 202.125 17.395 202.195 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 198.205 17.395 198.275 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 194.285 17.395 194.355 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 190.365 17.395 190.435 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 186.445 17.395 186.515 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 182.525 17.395 182.595 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 178.605 17.395 178.675 ;
        END
    END p377
    PIN p378
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 174.685 17.395 174.755 ;
        END
    END p378
    PIN p379
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 170.765 17.395 170.835 ;
        END
    END p379
    PIN p380
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 166.845 17.395 166.915 ;
        END
    END p380
    PIN p381
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 162.925 17.395 162.995 ;
        END
    END p381
    PIN p382
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 139.965 17.395 140.035 ;
        END
    END p382
    PIN p383
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 136.045 17.395 136.115 ;
        END
    END p383
    PIN p384
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 132.125 17.395 132.195 ;
        END
    END p384
    PIN p385
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 6.125 17.955 6.195 ;
        END
    END p385
    PIN p386
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 128.205 17.395 128.275 ;
        END
    END p386
    PIN p387
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 2.205 17.955 2.275 ;
        END
    END p387
    PIN p388
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 124.285 17.395 124.355 ;
        END
    END p388
    PIN p389
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 120.365 17.395 120.435 ;
        END
    END p389
    PIN p390
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 116.445 17.395 116.515 ;
        END
    END p390
    PIN p391
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 112.525 17.395 112.595 ;
        END
    END p391
    PIN p392
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 108.605 17.395 108.675 ;
        END
    END p392
    PIN p393
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 104.685 17.395 104.755 ;
        END
    END p393
    PIN p394
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 100.765 17.395 100.835 ;
        END
    END p394
    PIN p395
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 96.845 17.395 96.915 ;
        END
    END p395
    PIN p396
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 92.925 17.395 92.995 ;
        END
    END p396
    PIN p397
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 222.285 17.955 222.355 ;
        END
    END p397
    PIN p398
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 89.005 17.395 89.075 ;
        END
    END p398
    PIN p399
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 218.365 17.955 218.435 ;
        END
    END p399
    PIN p400
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 214.445 17.955 214.515 ;
        END
    END p400
    PIN p401
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 210.525 17.955 210.595 ;
        END
    END p401
    PIN p402
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 206.605 17.955 206.675 ;
        END
    END p402
    PIN p403
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 202.685 17.955 202.755 ;
        END
    END p403
    PIN p404
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 198.765 17.955 198.835 ;
        END
    END p404
    PIN p405
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 194.845 17.955 194.915 ;
        END
    END p405
    PIN p406
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 190.925 17.955 190.995 ;
        END
    END p406
    PIN p407
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 187.005 17.955 187.075 ;
        END
    END p407
    PIN p408
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 261.485 17.955 261.555 ;
        END
    END p408
    PIN p409
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 257.565 17.955 257.635 ;
        END
    END p409
    PIN p410
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 253.645 17.955 253.715 ;
        END
    END p410
    PIN p411
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 249.725 17.955 249.795 ;
        END
    END p411
    PIN p412
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 245.805 17.955 245.875 ;
        END
    END p412
    PIN p413
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 241.885 17.955 241.955 ;
        END
    END p413
    PIN p414
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 237.965 17.955 238.035 ;
        END
    END p414
    PIN p415
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 234.045 17.955 234.115 ;
        END
    END p415
    PIN p416
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 230.125 17.955 230.195 ;
        END
    END p416
    PIN p417
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 226.205 17.955 226.275 ;
        END
    END p417
    PIN p418
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 123.725 17.955 123.795 ;
        END
    END p418
    PIN p419
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 119.805 17.955 119.875 ;
        END
    END p419
    PIN p420
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 115.885 17.955 115.955 ;
        END
    END p420
    PIN p421
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 111.965 17.955 112.035 ;
        END
    END p421
    PIN p422
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 108.045 17.955 108.115 ;
        END
    END p422
    PIN p423
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 104.125 17.955 104.195 ;
        END
    END p423
    PIN p424
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 100.205 17.955 100.275 ;
        END
    END p424
    PIN p425
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 96.285 17.955 96.355 ;
        END
    END p425
    PIN p426
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 300.685 17.955 300.755 ;
        END
    END p426
    PIN p427
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 92.365 17.955 92.435 ;
        END
    END p427
    PIN p428
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 296.765 17.955 296.835 ;
        END
    END p428
    PIN p429
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 88.445 17.955 88.515 ;
        END
    END p429
    PIN p430
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 292.845 17.955 292.915 ;
        END
    END p430
    PIN p431
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 288.925 17.955 288.995 ;
        END
    END p431
    PIN p432
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 285.005 17.955 285.075 ;
        END
    END p432
    PIN p433
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 281.085 17.955 281.155 ;
        END
    END p433
    PIN p434
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 277.165 17.955 277.235 ;
        END
    END p434
    PIN p435
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 273.245 17.955 273.315 ;
        END
    END p435
    PIN p436
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 269.325 17.955 269.395 ;
        END
    END p436
    PIN p437
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 183.085 17.955 183.155 ;
        END
    END p437
    PIN p438
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 265.405 17.955 265.475 ;
        END
    END p438
    PIN p439
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 179.165 17.955 179.235 ;
        END
    END p439
    PIN p440
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 175.245 17.955 175.315 ;
        END
    END p440
    PIN p441
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 171.325 17.955 171.395 ;
        END
    END p441
    PIN p442
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 167.405 17.955 167.475 ;
        END
    END p442
    PIN p443
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 163.485 17.955 163.555 ;
        END
    END p443
    PIN p444
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 139.405 17.955 139.475 ;
        END
    END p444
    PIN p445
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 135.485 17.955 135.555 ;
        END
    END p445
    PIN p446
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 131.565 17.955 131.635 ;
        END
    END p446
    PIN p447
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 127.645 17.955 127.715 ;
        END
    END p447
    OBS
      LAYER via2 ;
        RECT  0 0 19.6 304.08 ;
      LAYER metal2 ;
        RECT  0 0 19.6 304.08 ;
      LAYER via1 ;
        RECT  0 0 19.6 304.08 ;
      LAYER metal1 ;
        RECT  0 0 19.6 304.08 ;
    END
END fake_macro_adaptec1_o211416

MACRO fake_macro_adaptec1_o211417
    CLASS BLOCK ;
    SIZE 15.12 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.805 0.595 252.875 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.205 0.595 233.275 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.325 0.595 178.395 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.725 0.595 158.795 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.085 0.595 141.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.485 0.595 121.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.965 13.475 154.035 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.685 13.475 153.755 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 152.005 13.475 152.075 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 142.205 13.475 142.275 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.925 13.475 169.995 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 154.245 14.035 154.315 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 295.085 13.475 295.155 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 291.165 13.475 291.235 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 287.245 13.475 287.315 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 283.325 13.475 283.395 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 279.405 13.475 279.475 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 275.485 13.475 275.555 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 271.565 13.475 271.635 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 267.645 13.475 267.715 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 263.725 13.475 263.795 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 259.805 13.475 259.875 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 85.085 13.475 85.155 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.165 13.475 81.235 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 77.245 13.475 77.315 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.325 13.475 73.395 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 69.405 13.475 69.475 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 65.485 13.475 65.555 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 61.565 13.475 61.635 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 57.645 13.475 57.715 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 53.725 13.475 53.795 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 49.805 13.475 49.875 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 45.885 13.475 45.955 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 41.965 13.475 42.035 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 38.045 13.475 38.115 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 34.125 13.475 34.195 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 30.205 13.475 30.275 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.285 13.475 26.355 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 22.365 13.475 22.435 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 18.445 13.475 18.515 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 14.525 13.475 14.595 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 10.605 13.475 10.675 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 6.685 13.475 6.755 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 2.765 13.475 2.835 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 255.885 13.475 255.955 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 251.965 13.475 252.035 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 248.045 13.475 248.115 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 244.125 13.475 244.195 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 240.205 13.475 240.275 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 236.285 13.475 236.355 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 232.365 13.475 232.435 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 228.445 13.475 228.515 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 224.525 13.475 224.595 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 220.605 13.475 220.675 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 216.685 13.475 216.755 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 212.765 13.475 212.835 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 208.845 13.475 208.915 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 204.925 13.475 204.995 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 201.005 13.475 201.075 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 197.085 13.475 197.155 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 193.165 13.475 193.235 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 189.245 13.475 189.315 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 185.325 13.475 185.395 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 181.405 13.475 181.475 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 177.485 13.475 177.555 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 173.565 13.475 173.635 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.645 13.475 169.715 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 165.725 13.475 165.795 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 161.805 13.475 161.875 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 157.885 13.475 157.955 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 139.965 13.475 140.035 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 136.045 13.475 136.115 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 132.125 13.475 132.195 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 128.205 13.475 128.275 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 124.285 13.475 124.355 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 120.365 13.475 120.435 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 116.445 13.475 116.515 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 112.525 13.475 112.595 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 108.605 13.475 108.675 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 104.685 13.475 104.755 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 100.765 13.475 100.835 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 96.845 13.475 96.915 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 92.925 13.475 92.995 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 89.005 13.475 89.075 ;
        END
    END p371
    OBS
      LAYER via2 ;
        RECT  0 0 15.12 299.04 ;
      LAYER metal2 ;
        RECT  0 0 15.12 299.04 ;
      LAYER via1 ;
        RECT  0 0 15.12 299.04 ;
      LAYER metal1 ;
        RECT  0 0 15.12 299.04 ;
    END
END fake_macro_adaptec1_o211417

MACRO fake_macro_adaptec1_o211418
    CLASS BLOCK ;
    SIZE 19.6 BY 304.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 158.165 17.395 158.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 300.685 0.595 300.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 157.045 17.395 157.115 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 156.765 0.595 156.835 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 156.205 0.595 156.275 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 159.845 0.595 159.915 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.405 0.595 160.475 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 142.205 17.395 142.275 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 169.925 17.395 169.995 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 145.005 0.595 145.075 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.845 0.595 271.915 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.765 0.595 275.835 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 285.285 0.595 285.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 281.365 0.595 281.435 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.165 0.595 137.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.925 0.595 267.995 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 265.685 0.595 265.755 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 246.085 0.595 246.155 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.325 0.595 234.395 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.885 0.595 220.955 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 199.045 0.595 199.115 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.605 0.595 185.675 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.085 0.595 162.155 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.725 0.595 228.795 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.805 0.595 224.875 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.645 0.595 218.715 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.045 0.595 213.115 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.125 0.595 209.195 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.685 0.595 181.755 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 179.445 0.595 179.515 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.845 0.595 173.915 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.685 0.595 167.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.445 0.595 291.515 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.245 0.595 252.315 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 238.245 0.595 238.315 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.205 0.595 205.275 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.605 0.595 171.675 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.285 0.595 201.355 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.445 0.595 193.515 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 191.205 0.595 191.275 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.285 0.595 299.355 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.365 0.595 295.435 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.525 0.595 287.595 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.085 0.595 260.155 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.165 0.595 256.235 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.325 0.595 248.395 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.485 0.595 240.555 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 163.485 0.595 163.555 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.405 0.595 167.475 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.325 0.595 171.395 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 175.245 0.595 175.315 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 179.165 0.595 179.235 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 183.085 0.595 183.155 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 187.005 0.595 187.075 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.925 0.595 190.995 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.845 0.595 194.915 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 198.765 0.595 198.835 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.685 0.595 202.755 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 206.605 0.595 206.675 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 210.525 0.595 210.595 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 214.445 0.595 214.515 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.365 0.595 218.435 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 222.285 0.595 222.355 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 226.205 0.595 226.275 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 230.125 0.595 230.195 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.045 0.595 234.115 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 237.965 0.595 238.035 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.885 0.595 241.955 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 245.805 0.595 245.875 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 249.725 0.595 249.795 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 253.645 0.595 253.715 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 257.565 0.595 257.635 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 261.485 0.595 261.555 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 265.405 0.595 265.475 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 269.325 0.595 269.395 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 273.245 0.595 273.315 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 277.165 0.595 277.235 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 281.085 0.595 281.155 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 285.005 0.595 285.075 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.925 0.595 288.995 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.845 0.595 292.915 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 296.765 0.595 296.835 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.565 0.595 299.635 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 152.285 17.395 152.355 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.445 0.595 151.515 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 150.885 0.595 150.955 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 152.285 0.595 152.355 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 159.005 16.275 159.075 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 186.725 16.275 186.795 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.925 0.595 162.995 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.845 0.595 166.915 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.765 0.595 170.835 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.685 0.595 174.755 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.605 0.595 178.675 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.525 0.595 182.595 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.445 0.595 186.515 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.365 0.595 190.435 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.285 0.595 194.355 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 198.205 0.595 198.275 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.125 0.595 202.195 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 206.045 0.595 206.115 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.965 0.595 210.035 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.885 0.595 213.955 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.805 0.595 217.875 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.725 0.595 221.795 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.645 0.595 225.715 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.565 0.595 229.635 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.485 0.595 233.555 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 237.405 0.595 237.475 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.325 0.595 241.395 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 245.245 0.595 245.315 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 249.165 0.595 249.235 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 253.085 0.595 253.155 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 257.005 0.595 257.075 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.925 0.595 260.995 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.845 0.595 264.915 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.765 0.595 268.835 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.365 0.595 288.435 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.685 0.595 272.755 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.285 0.595 292.355 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.605 0.595 276.675 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 296.205 0.595 296.275 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.525 0.595 280.595 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 300.125 0.595 300.195 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.445 0.595 284.515 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 265.405 17.955 265.475 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 85.085 17.395 85.155 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 81.165 17.395 81.235 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 77.245 17.395 77.315 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 73.325 17.395 73.395 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 69.405 17.395 69.475 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 65.485 17.395 65.555 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 61.565 17.395 61.635 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 57.645 17.395 57.715 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 53.725 17.395 53.795 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 49.805 17.395 49.875 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 45.885 17.395 45.955 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 41.965 17.395 42.035 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 38.045 17.395 38.115 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 34.125 17.395 34.195 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 30.205 17.395 30.275 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 26.285 17.395 26.355 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 22.365 17.395 22.435 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 18.445 17.395 18.515 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 14.525 17.395 14.595 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 10.605 17.395 10.675 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 6.685 17.395 6.755 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 2.765 17.395 2.835 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 300.125 17.395 300.195 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 296.205 17.395 296.275 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 292.285 17.395 292.355 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 288.365 17.395 288.435 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 284.445 17.395 284.515 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 280.525 17.395 280.595 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 276.605 17.395 276.675 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 272.685 17.395 272.755 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 268.765 17.395 268.835 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 264.845 17.395 264.915 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 45.325 17.955 45.395 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 41.405 17.955 41.475 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 37.485 17.955 37.555 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 33.565 17.955 33.635 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 29.645 17.955 29.715 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 25.725 17.955 25.795 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 21.805 17.955 21.875 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 17.885 17.955 17.955 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 13.965 17.955 14.035 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 10.045 17.955 10.115 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 260.925 17.395 260.995 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 257.005 17.395 257.075 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 253.085 17.395 253.155 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 249.165 17.395 249.235 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 245.245 17.395 245.315 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 241.325 17.395 241.395 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 237.405 17.395 237.475 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 84.525 17.955 84.595 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 233.485 17.395 233.555 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 80.605 17.955 80.675 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 229.565 17.395 229.635 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 76.685 17.955 76.755 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 225.645 17.395 225.715 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 72.765 17.955 72.835 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 68.845 17.955 68.915 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 64.925 17.955 64.995 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 61.005 17.955 61.075 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 57.085 17.955 57.155 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 53.165 17.955 53.235 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 49.245 17.955 49.315 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 221.725 17.395 221.795 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 217.805 17.395 217.875 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 213.885 17.395 213.955 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 209.965 17.395 210.035 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 206.045 17.395 206.115 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 202.125 17.395 202.195 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 198.205 17.395 198.275 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 194.285 17.395 194.355 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 190.365 17.395 190.435 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 186.445 17.395 186.515 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 182.525 17.395 182.595 ;
        END
    END p377
    PIN p378
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 178.605 17.395 178.675 ;
        END
    END p378
    PIN p379
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 174.685 17.395 174.755 ;
        END
    END p379
    PIN p380
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 170.765 17.395 170.835 ;
        END
    END p380
    PIN p381
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 166.845 17.395 166.915 ;
        END
    END p381
    PIN p382
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 162.925 17.395 162.995 ;
        END
    END p382
    PIN p383
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 139.965 17.395 140.035 ;
        END
    END p383
    PIN p384
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 6.125 17.955 6.195 ;
        END
    END p384
    PIN p385
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 136.045 17.395 136.115 ;
        END
    END p385
    PIN p386
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 2.205 17.955 2.275 ;
        END
    END p386
    PIN p387
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 132.125 17.395 132.195 ;
        END
    END p387
    PIN p388
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 128.205 17.395 128.275 ;
        END
    END p388
    PIN p389
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 124.285 17.395 124.355 ;
        END
    END p389
    PIN p390
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 120.365 17.395 120.435 ;
        END
    END p390
    PIN p391
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 116.445 17.395 116.515 ;
        END
    END p391
    PIN p392
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 112.525 17.395 112.595 ;
        END
    END p392
    PIN p393
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 108.605 17.395 108.675 ;
        END
    END p393
    PIN p394
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 104.685 17.395 104.755 ;
        END
    END p394
    PIN p395
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 100.765 17.395 100.835 ;
        END
    END p395
    PIN p396
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 222.285 17.955 222.355 ;
        END
    END p396
    PIN p397
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 96.845 17.395 96.915 ;
        END
    END p397
    PIN p398
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 218.365 17.955 218.435 ;
        END
    END p398
    PIN p399
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 92.925 17.395 92.995 ;
        END
    END p399
    PIN p400
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 214.445 17.955 214.515 ;
        END
    END p400
    PIN p401
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 89.005 17.395 89.075 ;
        END
    END p401
    PIN p402
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 210.525 17.955 210.595 ;
        END
    END p402
    PIN p403
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 206.605 17.955 206.675 ;
        END
    END p403
    PIN p404
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 202.685 17.955 202.755 ;
        END
    END p404
    PIN p405
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 198.765 17.955 198.835 ;
        END
    END p405
    PIN p406
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 194.845 17.955 194.915 ;
        END
    END p406
    PIN p407
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 190.925 17.955 190.995 ;
        END
    END p407
    PIN p408
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 187.005 17.955 187.075 ;
        END
    END p408
    PIN p409
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 261.485 17.955 261.555 ;
        END
    END p409
    PIN p410
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 257.565 17.955 257.635 ;
        END
    END p410
    PIN p411
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 253.645 17.955 253.715 ;
        END
    END p411
    PIN p412
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 249.725 17.955 249.795 ;
        END
    END p412
    PIN p413
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 245.805 17.955 245.875 ;
        END
    END p413
    PIN p414
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 241.885 17.955 241.955 ;
        END
    END p414
    PIN p415
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 237.965 17.955 238.035 ;
        END
    END p415
    PIN p416
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 234.045 17.955 234.115 ;
        END
    END p416
    PIN p417
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 230.125 17.955 230.195 ;
        END
    END p417
    PIN p418
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 226.205 17.955 226.275 ;
        END
    END p418
    PIN p419
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 123.725 17.955 123.795 ;
        END
    END p419
    PIN p420
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 119.805 17.955 119.875 ;
        END
    END p420
    PIN p421
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 115.885 17.955 115.955 ;
        END
    END p421
    PIN p422
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 111.965 17.955 112.035 ;
        END
    END p422
    PIN p423
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 108.045 17.955 108.115 ;
        END
    END p423
    PIN p424
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 104.125 17.955 104.195 ;
        END
    END p424
    PIN p425
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 100.205 17.955 100.275 ;
        END
    END p425
    PIN p426
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 96.285 17.955 96.355 ;
        END
    END p426
    PIN p427
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 92.365 17.955 92.435 ;
        END
    END p427
    PIN p428
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 88.445 17.955 88.515 ;
        END
    END p428
    PIN p429
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 183.085 17.955 183.155 ;
        END
    END p429
    PIN p430
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 179.165 17.955 179.235 ;
        END
    END p430
    PIN p431
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 175.245 17.955 175.315 ;
        END
    END p431
    PIN p432
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 171.325 17.955 171.395 ;
        END
    END p432
    PIN p433
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 167.405 17.955 167.475 ;
        END
    END p433
    PIN p434
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 163.485 17.955 163.555 ;
        END
    END p434
    PIN p435
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 139.405 17.955 139.475 ;
        END
    END p435
    PIN p436
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 135.485 17.955 135.555 ;
        END
    END p436
    PIN p437
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 131.565 17.955 131.635 ;
        END
    END p437
    PIN p438
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 300.685 17.955 300.755 ;
        END
    END p438
    PIN p439
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 127.645 17.955 127.715 ;
        END
    END p439
    PIN p440
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 296.765 17.955 296.835 ;
        END
    END p440
    PIN p441
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 292.845 17.955 292.915 ;
        END
    END p441
    PIN p442
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 288.925 17.955 288.995 ;
        END
    END p442
    PIN p443
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 285.005 17.955 285.075 ;
        END
    END p443
    PIN p444
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 281.085 17.955 281.155 ;
        END
    END p444
    PIN p445
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 277.165 17.955 277.235 ;
        END
    END p445
    PIN p446
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 273.245 17.955 273.315 ;
        END
    END p446
    PIN p447
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 269.325 17.955 269.395 ;
        END
    END p447
    OBS
      LAYER via2 ;
        RECT  0 0 19.6 304.08 ;
      LAYER metal2 ;
        RECT  0 0 19.6 304.08 ;
      LAYER via1 ;
        RECT  0 0 19.6 304.08 ;
      LAYER metal1 ;
        RECT  0 0 19.6 304.08 ;
    END
END fake_macro_adaptec1_o211418

MACRO fake_macro_adaptec1_o211419
    CLASS BLOCK ;
    SIZE 15.12 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.805 0.595 252.875 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.205 0.595 233.275 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.325 0.595 178.395 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.725 0.595 158.795 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.085 0.595 141.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.485 0.595 121.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.965 13.475 154.035 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.685 13.475 153.755 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 152.005 13.475 152.075 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 181.685 13.475 181.755 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 142.205 13.475 142.275 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.405 13.475 153.475 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 295.085 13.475 295.155 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 291.165 13.475 291.235 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 287.245 13.475 287.315 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 283.325 13.475 283.395 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 279.405 13.475 279.475 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 275.485 13.475 275.555 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 271.565 13.475 271.635 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 267.645 13.475 267.715 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 263.725 13.475 263.795 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 259.805 13.475 259.875 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 85.085 13.475 85.155 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.165 13.475 81.235 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 77.245 13.475 77.315 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.325 13.475 73.395 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 69.405 13.475 69.475 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 65.485 13.475 65.555 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 61.565 13.475 61.635 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 57.645 13.475 57.715 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 53.725 13.475 53.795 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 49.805 13.475 49.875 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 45.885 13.475 45.955 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 41.965 13.475 42.035 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 38.045 13.475 38.115 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 34.125 13.475 34.195 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 30.205 13.475 30.275 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.285 13.475 26.355 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 22.365 13.475 22.435 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 18.445 13.475 18.515 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 14.525 13.475 14.595 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 10.605 13.475 10.675 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 6.685 13.475 6.755 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 2.765 13.475 2.835 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 255.885 13.475 255.955 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 251.965 13.475 252.035 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 248.045 13.475 248.115 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 244.125 13.475 244.195 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 240.205 13.475 240.275 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 236.285 13.475 236.355 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 232.365 13.475 232.435 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 228.445 13.475 228.515 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 224.525 13.475 224.595 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 220.605 13.475 220.675 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 216.685 13.475 216.755 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 212.765 13.475 212.835 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 208.845 13.475 208.915 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 204.925 13.475 204.995 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 201.005 13.475 201.075 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 197.085 13.475 197.155 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 193.165 13.475 193.235 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 189.245 13.475 189.315 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 185.325 13.475 185.395 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 181.405 13.475 181.475 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 177.485 13.475 177.555 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 173.565 13.475 173.635 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.645 13.475 169.715 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 165.725 13.475 165.795 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 161.805 13.475 161.875 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 157.885 13.475 157.955 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 139.965 13.475 140.035 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 136.045 13.475 136.115 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 132.125 13.475 132.195 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 128.205 13.475 128.275 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 124.285 13.475 124.355 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 120.365 13.475 120.435 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 116.445 13.475 116.515 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 112.525 13.475 112.595 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 108.605 13.475 108.675 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 104.685 13.475 104.755 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 100.765 13.475 100.835 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 96.845 13.475 96.915 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 92.925 13.475 92.995 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 89.005 13.475 89.075 ;
        END
    END p371
    OBS
      LAYER via2 ;
        RECT  0 0 15.12 299.04 ;
      LAYER metal2 ;
        RECT  0 0 15.12 299.04 ;
      LAYER via1 ;
        RECT  0 0 15.12 299.04 ;
      LAYER metal1 ;
        RECT  0 0 15.12 299.04 ;
    END
END fake_macro_adaptec1_o211419

MACRO fake_macro_adaptec1_o211420
    CLASS BLOCK ;
    SIZE 19.6 BY 304.08 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 158.165 17.395 158.235 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 300.685 0.595 300.755 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 159.005 16.275 159.075 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 157.045 17.395 157.115 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 156.765 0.595 156.835 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 156.205 0.595 156.275 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 159.845 0.595 159.915 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 142.205 17.395 142.275 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 169.925 17.395 169.995 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 145.005 0.595 145.075 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.765 0.595 275.835 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 48.965 0.595 49.035 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 281.365 0.595 281.435 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.845 0.595 271.915 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.325 0.595 248.395 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.885 0.595 220.955 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 199.045 0.595 199.115 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 179.445 0.595 179.515 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.525 0.595 287.595 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.165 0.595 256.235 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.725 0.595 228.795 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.205 0.595 205.275 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.605 0.595 185.675 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.085 0.595 162.155 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.165 0.595 137.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.805 0.595 224.875 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.645 0.595 218.715 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.045 0.595 213.115 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.125 0.595 209.195 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.285 0.595 201.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.445 0.595 193.515 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 191.205 0.595 191.275 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.685 0.595 181.755 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.845 0.595 173.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.605 0.595 171.675 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.685 0.595 167.755 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.285 0.595 299.355 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.365 0.595 295.435 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.445 0.595 291.515 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.925 0.595 267.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 265.685 0.595 265.755 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.085 0.595 260.155 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.245 0.595 252.315 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 246.085 0.595 246.155 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.485 0.595 240.555 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 238.245 0.595 238.315 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.325 0.595 234.395 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 152.285 17.395 152.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.445 0.595 151.515 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 150.885 0.595 150.955 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 152.285 0.595 152.355 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  16.205 186.725 16.275 186.795 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.925 0.595 162.995 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.845 0.595 166.915 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.765 0.595 170.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.685 0.595 174.755 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.605 0.595 178.675 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.525 0.595 182.595 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.445 0.595 186.515 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.365 0.595 190.435 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.285 0.595 194.355 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 198.205 0.595 198.275 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.125 0.595 202.195 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 206.045 0.595 206.115 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.965 0.595 210.035 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.885 0.595 213.955 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.805 0.595 217.875 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.725 0.595 221.795 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.645 0.595 225.715 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.565 0.595 229.635 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.485 0.595 233.555 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 237.405 0.595 237.475 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.325 0.595 241.395 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 245.245 0.595 245.315 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 249.165 0.595 249.235 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 253.085 0.595 253.155 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 257.005 0.595 257.075 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.925 0.595 260.995 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.845 0.595 264.915 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.765 0.595 268.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.365 0.595 288.435 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.685 0.595 272.755 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.285 0.595 292.355 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.605 0.595 276.675 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 296.205 0.595 296.275 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.525 0.595 280.595 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 300.125 0.595 300.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.445 0.595 284.515 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.405 0.595 160.475 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 285.285 0.595 285.355 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.685 0.595 111.755 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 163.485 0.595 163.555 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 167.405 0.595 167.475 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 171.325 0.595 171.395 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 175.245 0.595 175.315 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 179.165 0.595 179.235 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 183.085 0.595 183.155 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 187.005 0.595 187.075 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.925 0.595 190.995 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.845 0.595 194.915 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 198.765 0.595 198.835 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 202.685 0.595 202.755 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 206.605 0.595 206.675 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 210.525 0.595 210.595 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 214.445 0.595 214.515 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 218.365 0.595 218.435 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 222.285 0.595 222.355 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 226.205 0.595 226.275 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 230.125 0.595 230.195 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 234.045 0.595 234.115 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 237.965 0.595 238.035 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.885 0.595 241.955 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 245.805 0.595 245.875 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 249.725 0.595 249.795 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 253.645 0.595 253.715 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 257.565 0.595 257.635 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 261.485 0.595 261.555 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p285
    PIN p286
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 265.405 0.595 265.475 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p287
    PIN p288
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 269.325 0.595 269.395 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p289
    PIN p290
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 273.245 0.595 273.315 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p291
    PIN p292
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 277.165 0.595 277.235 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p293
    PIN p294
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 281.085 0.595 281.155 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p295
    PIN p296
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 285.005 0.595 285.075 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.925 0.595 288.995 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.845 0.595 292.915 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 296.765 0.595 296.835 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 299.565 0.595 299.635 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 85.085 17.395 85.155 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 81.165 17.395 81.235 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 77.245 17.395 77.315 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 73.325 17.395 73.395 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 69.405 17.395 69.475 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 65.485 17.395 65.555 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 61.565 17.395 61.635 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 57.645 17.395 57.715 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 53.725 17.395 53.795 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 49.805 17.395 49.875 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 45.885 17.395 45.955 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 41.965 17.395 42.035 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 38.045 17.395 38.115 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 34.125 17.395 34.195 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 30.205 17.395 30.275 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 26.285 17.395 26.355 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 22.365 17.395 22.435 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 18.445 17.395 18.515 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 14.525 17.395 14.595 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 10.605 17.395 10.675 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 6.685 17.395 6.755 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 2.765 17.395 2.835 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 45.325 17.955 45.395 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 41.405 17.955 41.475 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 37.485 17.955 37.555 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 33.565 17.955 33.635 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 29.645 17.955 29.715 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 300.125 17.395 300.195 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 25.725 17.955 25.795 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 296.205 17.395 296.275 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 21.805 17.955 21.875 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 292.285 17.395 292.355 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 17.885 17.955 17.955 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 260.925 17.395 260.995 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 288.365 17.395 288.435 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 13.965 17.955 14.035 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 257.005 17.395 257.075 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 284.445 17.395 284.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 10.045 17.955 10.115 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 253.085 17.395 253.155 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 280.525 17.395 280.595 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 249.165 17.395 249.235 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 276.605 17.395 276.675 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 245.245 17.395 245.315 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 272.685 17.395 272.755 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 241.325 17.395 241.395 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 268.765 17.395 268.835 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 237.405 17.395 237.475 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 264.845 17.395 264.915 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 233.485 17.395 233.555 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 229.565 17.395 229.635 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 84.525 17.955 84.595 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 225.645 17.395 225.715 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 80.605 17.955 80.675 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 76.685 17.955 76.755 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 72.765 17.955 72.835 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 68.845 17.955 68.915 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 64.925 17.955 64.995 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 61.005 17.955 61.075 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 57.085 17.955 57.155 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 221.725 17.395 221.795 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 53.165 17.955 53.235 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 217.805 17.395 217.875 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 49.245 17.955 49.315 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 213.885 17.395 213.955 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 209.965 17.395 210.035 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 206.045 17.395 206.115 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 202.125 17.395 202.195 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 198.205 17.395 198.275 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 194.285 17.395 194.355 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 190.365 17.395 190.435 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 186.445 17.395 186.515 ;
        END
    END p375
    PIN p376
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 182.525 17.395 182.595 ;
        END
    END p376
    PIN p377
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 178.605 17.395 178.675 ;
        END
    END p377
    PIN p378
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 174.685 17.395 174.755 ;
        END
    END p378
    PIN p379
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 170.765 17.395 170.835 ;
        END
    END p379
    PIN p380
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 166.845 17.395 166.915 ;
        END
    END p380
    PIN p381
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 162.925 17.395 162.995 ;
        END
    END p381
    PIN p382
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 139.965 17.395 140.035 ;
        END
    END p382
    PIN p383
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 136.045 17.395 136.115 ;
        END
    END p383
    PIN p384
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 132.125 17.395 132.195 ;
        END
    END p384
    PIN p385
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 6.125 17.955 6.195 ;
        END
    END p385
    PIN p386
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 128.205 17.395 128.275 ;
        END
    END p386
    PIN p387
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 2.205 17.955 2.275 ;
        END
    END p387
    PIN p388
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 124.285 17.395 124.355 ;
        END
    END p388
    PIN p389
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 120.365 17.395 120.435 ;
        END
    END p389
    PIN p390
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 116.445 17.395 116.515 ;
        END
    END p390
    PIN p391
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 112.525 17.395 112.595 ;
        END
    END p391
    PIN p392
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 108.605 17.395 108.675 ;
        END
    END p392
    PIN p393
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 104.685 17.395 104.755 ;
        END
    END p393
    PIN p394
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 100.765 17.395 100.835 ;
        END
    END p394
    PIN p395
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 96.845 17.395 96.915 ;
        END
    END p395
    PIN p396
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 92.925 17.395 92.995 ;
        END
    END p396
    PIN p397
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 222.285 17.955 222.355 ;
        END
    END p397
    PIN p398
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.325 89.005 17.395 89.075 ;
        END
    END p398
    PIN p399
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 218.365 17.955 218.435 ;
        END
    END p399
    PIN p400
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 214.445 17.955 214.515 ;
        END
    END p400
    PIN p401
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 210.525 17.955 210.595 ;
        END
    END p401
    PIN p402
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 206.605 17.955 206.675 ;
        END
    END p402
    PIN p403
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 202.685 17.955 202.755 ;
        END
    END p403
    PIN p404
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 198.765 17.955 198.835 ;
        END
    END p404
    PIN p405
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 194.845 17.955 194.915 ;
        END
    END p405
    PIN p406
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 190.925 17.955 190.995 ;
        END
    END p406
    PIN p407
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 187.005 17.955 187.075 ;
        END
    END p407
    PIN p408
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 261.485 17.955 261.555 ;
        END
    END p408
    PIN p409
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 257.565 17.955 257.635 ;
        END
    END p409
    PIN p410
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 253.645 17.955 253.715 ;
        END
    END p410
    PIN p411
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 249.725 17.955 249.795 ;
        END
    END p411
    PIN p412
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 245.805 17.955 245.875 ;
        END
    END p412
    PIN p413
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 241.885 17.955 241.955 ;
        END
    END p413
    PIN p414
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 237.965 17.955 238.035 ;
        END
    END p414
    PIN p415
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 234.045 17.955 234.115 ;
        END
    END p415
    PIN p416
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 230.125 17.955 230.195 ;
        END
    END p416
    PIN p417
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 226.205 17.955 226.275 ;
        END
    END p417
    PIN p418
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 123.725 17.955 123.795 ;
        END
    END p418
    PIN p419
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 119.805 17.955 119.875 ;
        END
    END p419
    PIN p420
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 115.885 17.955 115.955 ;
        END
    END p420
    PIN p421
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 111.965 17.955 112.035 ;
        END
    END p421
    PIN p422
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 108.045 17.955 108.115 ;
        END
    END p422
    PIN p423
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 104.125 17.955 104.195 ;
        END
    END p423
    PIN p424
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 100.205 17.955 100.275 ;
        END
    END p424
    PIN p425
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 96.285 17.955 96.355 ;
        END
    END p425
    PIN p426
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 300.685 17.955 300.755 ;
        END
    END p426
    PIN p427
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 92.365 17.955 92.435 ;
        END
    END p427
    PIN p428
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 296.765 17.955 296.835 ;
        END
    END p428
    PIN p429
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 88.445 17.955 88.515 ;
        END
    END p429
    PIN p430
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 292.845 17.955 292.915 ;
        END
    END p430
    PIN p431
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 288.925 17.955 288.995 ;
        END
    END p431
    PIN p432
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 285.005 17.955 285.075 ;
        END
    END p432
    PIN p433
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 281.085 17.955 281.155 ;
        END
    END p433
    PIN p434
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 277.165 17.955 277.235 ;
        END
    END p434
    PIN p435
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 273.245 17.955 273.315 ;
        END
    END p435
    PIN p436
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 269.325 17.955 269.395 ;
        END
    END p436
    PIN p437
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 183.085 17.955 183.155 ;
        END
    END p437
    PIN p438
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 265.405 17.955 265.475 ;
        END
    END p438
    PIN p439
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 179.165 17.955 179.235 ;
        END
    END p439
    PIN p440
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 175.245 17.955 175.315 ;
        END
    END p440
    PIN p441
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 171.325 17.955 171.395 ;
        END
    END p441
    PIN p442
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 167.405 17.955 167.475 ;
        END
    END p442
    PIN p443
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 163.485 17.955 163.555 ;
        END
    END p443
    PIN p444
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 139.405 17.955 139.475 ;
        END
    END p444
    PIN p445
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 135.485 17.955 135.555 ;
        END
    END p445
    PIN p446
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 131.565 17.955 131.635 ;
        END
    END p446
    PIN p447
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  17.885 127.645 17.955 127.715 ;
        END
    END p447
    OBS
      LAYER via2 ;
        RECT  0 0 19.6 304.08 ;
      LAYER metal2 ;
        RECT  0 0 19.6 304.08 ;
      LAYER via1 ;
        RECT  0 0 19.6 304.08 ;
      LAYER metal1 ;
        RECT  0 0 19.6 304.08 ;
    END
END fake_macro_adaptec1_o211420

MACRO fake_macro_adaptec1_o211421
    CLASS BLOCK ;
    SIZE 15.12 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.805 0.595 252.875 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.205 0.595 233.275 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.325 0.595 178.395 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.725 0.595 158.795 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.085 0.595 141.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.485 0.595 121.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.965 13.475 154.035 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 153.685 13.475 153.755 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 152.005 13.475 152.075 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 142.205 13.475 142.275 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.925 13.475 169.995 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.965 154.245 14.035 154.315 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 295.085 13.475 295.155 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 291.165 13.475 291.235 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 287.245 13.475 287.315 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 283.325 13.475 283.395 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 279.405 13.475 279.475 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 275.485 13.475 275.555 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 271.565 13.475 271.635 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 267.645 13.475 267.715 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 263.725 13.475 263.795 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 259.805 13.475 259.875 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 85.085 13.475 85.155 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 81.165 13.475 81.235 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 77.245 13.475 77.315 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 73.325 13.475 73.395 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 69.405 13.475 69.475 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 65.485 13.475 65.555 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 61.565 13.475 61.635 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 57.645 13.475 57.715 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 53.725 13.475 53.795 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 49.805 13.475 49.875 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 45.885 13.475 45.955 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 41.965 13.475 42.035 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 38.045 13.475 38.115 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 34.125 13.475 34.195 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 30.205 13.475 30.275 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 26.285 13.475 26.355 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 22.365 13.475 22.435 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 18.445 13.475 18.515 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 14.525 13.475 14.595 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 10.605 13.475 10.675 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 6.685 13.475 6.755 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 2.765 13.475 2.835 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 255.885 13.475 255.955 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 251.965 13.475 252.035 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 248.045 13.475 248.115 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 244.125 13.475 244.195 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 240.205 13.475 240.275 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 236.285 13.475 236.355 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 232.365 13.475 232.435 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 228.445 13.475 228.515 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 224.525 13.475 224.595 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 220.605 13.475 220.675 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 216.685 13.475 216.755 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 212.765 13.475 212.835 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 208.845 13.475 208.915 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 204.925 13.475 204.995 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 201.005 13.475 201.075 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 197.085 13.475 197.155 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 193.165 13.475 193.235 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 189.245 13.475 189.315 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 185.325 13.475 185.395 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 181.405 13.475 181.475 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 177.485 13.475 177.555 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 173.565 13.475 173.635 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 169.645 13.475 169.715 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 165.725 13.475 165.795 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 161.805 13.475 161.875 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 157.885 13.475 157.955 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 139.965 13.475 140.035 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 136.045 13.475 136.115 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 132.125 13.475 132.195 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 128.205 13.475 128.275 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 124.285 13.475 124.355 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 120.365 13.475 120.435 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 116.445 13.475 116.515 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 112.525 13.475 112.595 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 108.605 13.475 108.675 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 104.685 13.475 104.755 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 100.765 13.475 100.835 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 96.845 13.475 96.915 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 92.925 13.475 92.995 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  13.405 89.005 13.475 89.075 ;
        END
    END p371
    OBS
      LAYER via2 ;
        RECT  0 0 15.12 299.04 ;
      LAYER metal2 ;
        RECT  0 0 15.12 299.04 ;
      LAYER via1 ;
        RECT  0 0 15.12 299.04 ;
      LAYER metal1 ;
        RECT  0 0 15.12 299.04 ;
    END
END fake_macro_adaptec1_o211421

MACRO fake_macro_adaptec1_o211422
    CLASS BLOCK ;
    SIZE 11.2 BY 142.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.845 0.595 117.915 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.005 0.595 110.075 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.085 0.595 106.155 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.565 0.595 82.635 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.685 0.595 62.755 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 56.805 0.595 56.875 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.405 0.595 27.475 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 75.565 9.555 75.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 103.285 9.555 103.355 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 73.605 9.555 73.675 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 75.285 9.555 75.355 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.045 0.595 80.115 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.965 0.595 84.035 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.925 0.595 78.995 ;
        END
    END p73
    PIN p74
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.885 0.595 87.955 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.845 0.595 82.915 ;
        END
    END p75
    PIN p76
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.805 0.595 91.875 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.765 0.595 86.835 ;
        END
    END p77
    PIN p78
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.725 0.595 95.795 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.685 0.595 90.755 ;
        END
    END p79
    PIN p80
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.645 0.595 99.715 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.605 0.595 94.675 ;
        END
    END p81
    PIN p82
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.565 0.595 103.635 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 98.525 0.595 98.595 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.485 0.595 107.555 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 102.445 0.595 102.515 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.405 0.595 111.475 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.365 0.595 106.435 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.325 0.595 115.395 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.285 0.595 110.355 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.245 0.595 119.315 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.205 0.595 114.275 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.165 0.595 123.235 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.125 0.595 118.195 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.085 0.595 127.155 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.045 0.595 122.115 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.005 0.595 131.075 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.965 0.595 126.035 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.925 0.595 134.995 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.885 0.595 129.955 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.845 0.595 138.915 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.805 0.595 133.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.725 0.595 137.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 79.485 0.595 79.555 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.405 0.595 83.475 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.325 0.595 87.395 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.245 0.595 91.315 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.165 0.595 95.235 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.085 0.595 99.155 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.005 0.595 103.075 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.925 0.595 106.995 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.845 0.595 110.915 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.765 0.595 114.835 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.685 0.595 118.755 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.605 0.595 122.675 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.525 0.595 126.595 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.445 0.595 130.515 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.365 0.595 134.435 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.285 0.595 138.355 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 63.805 9.555 63.875 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 75.005 9.555 75.075 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 99.085 9.555 99.155 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 95.165 9.555 95.235 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 91.245 9.555 91.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 87.325 9.555 87.395 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 83.405 9.555 83.475 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 79.485 9.555 79.555 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 61.565 9.555 61.635 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 57.645 9.555 57.715 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 53.725 9.555 53.795 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 49.805 9.555 49.875 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 45.885 9.555 45.955 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 38.045 9.555 38.115 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 34.125 9.555 34.195 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 30.205 9.555 30.275 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 26.285 9.555 26.355 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 22.365 9.555 22.435 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 18.445 9.555 18.515 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 14.525 9.555 14.595 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.605 9.555 10.675 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 6.685 9.555 6.755 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.765 9.555 2.835 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.285 9.555 138.355 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 134.365 9.555 134.435 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 126.525 9.555 126.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 122.605 9.555 122.675 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 118.685 9.555 118.755 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 114.765 9.555 114.835 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 110.845 9.555 110.915 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 106.925 9.555 106.995 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 103.005 9.555 103.075 ;
        END
    END p169
    OBS
      LAYER via2 ;
        RECT  0 0 11.2 142.8 ;
      LAYER metal2 ;
        RECT  0 0 11.2 142.8 ;
      LAYER via1 ;
        RECT  0 0 11.2 142.8 ;
      LAYER metal1 ;
        RECT  0 0 11.2 142.8 ;
    END
END fake_macro_adaptec1_o211422

MACRO fake_macro_adaptec1_o211423
    CLASS BLOCK ;
    SIZE 71.4 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.125 69.475 153.195 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 153.965 68.915 154.035 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.005 69.475 152.075 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.085 69.475 148.155 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 149.485 3.395 149.555 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 150.605 2.275 150.675 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.245 2.275 119.315 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.405 2.275 111.475 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.565 2.275 103.635 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 95.725 2.275 95.795 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 87.885 2.275 87.955 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.045 2.275 80.115 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.205 2.275 72.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.365 2.275 64.435 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.685 2.275 195.755 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 187.845 2.275 187.915 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.005 2.275 180.075 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.165 2.275 172.235 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.325 2.275 164.395 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.485 2.275 156.555 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.925 2.275 134.995 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.085 2.275 127.155 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.405 2.275 258.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.565 2.275 250.635 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 242.725 2.275 242.795 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 234.885 2.275 234.955 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.045 2.275 227.115 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.205 2.275 219.275 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.365 2.275 211.435 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.525 2.275 203.595 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 289.765 2.275 289.835 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 281.925 2.275 281.995 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.085 2.275 274.155 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.245 2.275 266.315 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 181.685 68.915 181.755 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.605 1.155 3.675 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.445 1.155 11.515 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.285 1.155 19.355 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.125 1.155 27.195 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.965 1.155 35.035 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.805 1.155 42.875 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.645 1.155 50.715 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.485 1.155 58.555 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.325 1.155 66.395 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.165 1.155 74.235 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.005 1.155 82.075 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.845 1.155 89.915 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.525 1.155 105.595 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.365 1.155 113.435 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.205 1.155 121.275 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.045 1.155 129.115 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.485 1.155 184.555 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.165 1.155 200.235 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.525 1.155 231.595 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.165 0.595 144.235 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.205 68.915 142.275 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.365 3.955 148.435 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.245 2.275 147.315 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 181.405 70.035 181.475 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 173.565 70.035 173.635 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 164.605 70.035 164.675 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 157.885 70.035 157.955 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.965 70.035 140.035 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 132.125 70.035 132.195 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 124.285 70.035 124.355 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 116.445 70.035 116.515 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 108.605 70.035 108.675 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 100.765 70.035 100.835 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 94.045 70.035 94.115 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 85.085 70.035 85.155 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 77.245 70.035 77.315 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 70.525 70.035 70.595 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 61.565 70.035 61.635 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 53.725 70.035 53.795 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 47.005 70.035 47.075 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 38.045 70.035 38.115 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 30.205 70.035 30.275 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 23.485 70.035 23.555 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 14.525 70.035 14.595 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 6.685 70.035 6.755 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 291.165 70.035 291.235 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 283.325 70.035 283.395 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 275.485 70.035 275.555 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 267.645 70.035 267.715 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 259.805 70.035 259.875 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 251.965 70.035 252.035 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 244.125 70.035 244.195 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 235.165 70.035 235.235 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 228.445 70.035 228.515 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 220.605 70.035 220.675 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 211.645 70.035 211.715 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 204.925 70.035 204.995 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 197.085 70.035 197.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 188.125 70.035 188.195 ;
        END
    END p199
    OBS
      LAYER via2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER via1 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal1 ;
        RECT  0 0 71.54 299.04 ;
    END
END fake_macro_adaptec1_o211423

MACRO fake_macro_adaptec1_o211424
    CLASS BLOCK ;
    SIZE 71.4 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.125 69.475 153.195 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.005 69.475 152.075 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.085 69.475 148.155 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 149.485 3.395 149.555 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 150.605 2.275 150.675 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 234.885 2.275 234.955 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 242.725 2.275 242.795 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.565 2.275 250.635 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.405 2.275 258.475 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.245 2.275 266.315 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.165 0.595 144.235 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.205 68.915 142.275 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.365 3.955 148.435 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.245 2.275 147.315 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.085 2.275 274.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 87.885 2.275 87.955 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.045 2.275 80.115 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.205 2.275 72.275 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.365 2.275 64.435 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 281.925 2.275 281.995 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.325 2.275 164.395 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.485 2.275 156.555 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.925 2.275 134.995 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.085 2.275 127.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.245 2.275 119.315 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.405 2.275 111.475 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.565 2.275 103.635 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 95.725 2.275 95.795 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 289.765 2.275 289.835 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.045 2.275 227.115 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.205 2.275 219.275 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.365 2.275 211.435 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.525 2.275 203.595 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.685 2.275 195.755 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 187.845 2.275 187.915 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.005 2.275 180.075 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.165 2.275 172.235 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 153.965 68.915 154.035 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.605 1.155 3.675 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.445 1.155 11.515 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.285 1.155 19.355 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.125 1.155 27.195 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.965 1.155 35.035 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.805 1.155 42.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.645 1.155 50.715 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.485 1.155 58.555 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.325 1.155 66.395 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.165 1.155 74.235 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.005 1.155 82.075 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.845 1.155 89.915 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.525 1.155 105.595 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.365 1.155 113.435 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.205 1.155 121.275 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.045 1.155 129.115 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.485 1.155 184.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.165 1.155 200.235 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.525 1.155 231.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 181.685 68.915 181.755 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 291.165 70.035 291.235 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 283.325 70.035 283.395 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 275.485 70.035 275.555 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 267.645 70.035 267.715 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 259.805 70.035 259.875 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 251.965 70.035 252.035 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 244.125 70.035 244.195 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 235.165 70.035 235.235 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 228.445 70.035 228.515 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 220.605 70.035 220.675 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 211.645 70.035 211.715 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 204.925 70.035 204.995 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 197.085 70.035 197.155 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 188.125 70.035 188.195 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 181.405 70.035 181.475 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 173.565 70.035 173.635 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 164.605 70.035 164.675 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 157.885 70.035 157.955 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.965 70.035 140.035 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 132.125 70.035 132.195 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 124.285 70.035 124.355 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 116.445 70.035 116.515 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 108.605 70.035 108.675 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 100.765 70.035 100.835 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 94.045 70.035 94.115 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 85.085 70.035 85.155 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 77.245 70.035 77.315 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 70.525 70.035 70.595 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 61.565 70.035 61.635 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 53.725 70.035 53.795 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 47.005 70.035 47.075 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 38.045 70.035 38.115 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 30.205 70.035 30.275 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 23.485 70.035 23.555 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 14.525 70.035 14.595 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 6.685 70.035 6.755 ;
        END
    END p199
    OBS
      LAYER via2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER via1 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal1 ;
        RECT  0 0 71.54 299.04 ;
    END
END fake_macro_adaptec1_o211424

MACRO fake_macro_adaptec1_o211425
    CLASS BLOCK ;
    SIZE 71.4 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.005 69.475 152.075 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.085 69.475 148.155 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 149.485 3.395 149.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 150.605 2.275 150.675 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.605 1.155 3.675 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.445 1.155 11.515 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.285 1.155 19.355 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.125 1.155 27.195 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.965 1.155 35.035 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.805 1.155 42.875 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.645 1.155 50.715 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.485 1.155 58.555 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.325 1.155 66.395 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.165 1.155 74.235 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.005 1.155 82.075 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.845 1.155 89.915 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.525 1.155 105.595 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.365 1.155 113.435 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.205 1.155 121.275 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.045 1.155 129.115 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.485 1.155 184.555 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.165 1.155 200.235 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.525 1.155 231.595 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.165 0.595 144.235 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.205 68.915 142.275 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.365 3.955 148.435 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.245 2.275 147.315 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 153.965 68.915 154.035 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.245 2.275 119.315 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.405 2.275 111.475 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.565 2.275 103.635 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 95.725 2.275 95.795 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 87.885 2.275 87.955 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.045 2.275 80.115 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.205 2.275 72.275 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.365 2.275 64.435 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.685 2.275 195.755 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 187.845 2.275 187.915 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.005 2.275 180.075 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.165 2.275 172.235 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.325 2.275 164.395 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.485 2.275 156.555 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.925 2.275 134.995 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.085 2.275 127.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.405 2.275 258.475 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.565 2.275 250.635 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 242.725 2.275 242.795 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 234.885 2.275 234.955 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.045 2.275 227.115 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.205 2.275 219.275 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.365 2.275 211.435 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.525 2.275 203.595 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 289.765 2.275 289.835 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 281.925 2.275 281.995 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.085 2.275 274.155 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.245 2.275 266.315 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 181.685 68.915 181.755 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.125 69.475 153.195 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 181.405 70.035 181.475 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 173.565 70.035 173.635 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 164.605 70.035 164.675 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 157.885 70.035 157.955 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.965 70.035 140.035 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 132.125 70.035 132.195 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 124.285 70.035 124.355 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 116.445 70.035 116.515 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 108.605 70.035 108.675 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 100.765 70.035 100.835 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 94.045 70.035 94.115 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 85.085 70.035 85.155 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 77.245 70.035 77.315 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 70.525 70.035 70.595 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 61.565 70.035 61.635 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 53.725 70.035 53.795 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 47.005 70.035 47.075 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 38.045 70.035 38.115 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 30.205 70.035 30.275 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 23.485 70.035 23.555 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 14.525 70.035 14.595 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 6.685 70.035 6.755 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 291.165 70.035 291.235 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 283.325 70.035 283.395 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 275.485 70.035 275.555 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 267.645 70.035 267.715 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 259.805 70.035 259.875 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 251.965 70.035 252.035 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 244.125 70.035 244.195 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 235.165 70.035 235.235 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 228.445 70.035 228.515 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 220.605 70.035 220.675 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 211.645 70.035 211.715 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 204.925 70.035 204.995 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 197.085 70.035 197.155 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 188.125 70.035 188.195 ;
        END
    END p199
    OBS
      LAYER via2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER via1 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal1 ;
        RECT  0 0 71.54 299.04 ;
    END
END fake_macro_adaptec1_o211425

MACRO fake_macro_adaptec1_o211426
    CLASS BLOCK ;
    SIZE 71.4 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.005 69.475 152.075 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.085 69.475 148.155 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 149.485 3.395 149.555 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 150.605 2.275 150.675 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.165 0.595 144.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.205 68.915 142.275 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.365 3.955 148.435 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.245 2.275 147.315 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.605 1.155 3.675 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.445 1.155 11.515 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.285 1.155 19.355 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.125 1.155 27.195 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.965 1.155 35.035 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.805 1.155 42.875 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.645 1.155 50.715 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.485 1.155 58.555 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.325 1.155 66.395 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.165 1.155 74.235 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.005 1.155 82.075 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.845 1.155 89.915 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.365 1.155 113.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.045 1.155 129.115 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.485 1.155 184.555 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.165 1.155 200.235 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.525 1.155 231.595 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 153.965 68.915 154.035 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.245 2.275 266.315 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.085 2.275 274.155 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 87.885 2.275 87.955 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.045 2.275 80.115 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.205 2.275 72.275 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.365 2.275 64.435 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 281.925 2.275 281.995 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.325 2.275 164.395 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.485 2.275 156.555 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.925 2.275 134.995 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.085 2.275 127.155 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.245 2.275 119.315 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.405 2.275 111.475 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.565 2.275 103.635 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 95.725 2.275 95.795 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.045 2.275 227.115 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.205 2.275 219.275 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.365 2.275 211.435 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.525 2.275 203.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.685 2.275 195.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 187.845 2.275 187.915 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.005 2.275 180.075 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.165 2.275 172.235 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 234.885 2.275 234.955 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 242.725 2.275 242.795 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.565 2.275 250.635 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.405 2.275 258.475 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 289.765 2.275 289.835 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 181.685 68.915 181.755 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.525 1.155 105.595 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.205 1.155 121.275 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.125 69.475 153.195 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 211.645 70.035 211.715 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 204.925 70.035 204.995 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 197.085 70.035 197.155 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 188.125 70.035 188.195 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 181.405 70.035 181.475 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 173.565 70.035 173.635 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 164.605 70.035 164.675 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 157.885 70.035 157.955 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.965 70.035 140.035 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 132.125 70.035 132.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 124.285 70.035 124.355 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 116.445 70.035 116.515 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 108.605 70.035 108.675 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 100.765 70.035 100.835 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 94.045 70.035 94.115 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 85.085 70.035 85.155 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 77.245 70.035 77.315 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 70.525 70.035 70.595 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 61.565 70.035 61.635 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 53.725 70.035 53.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 47.005 70.035 47.075 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 38.045 70.035 38.115 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 30.205 70.035 30.275 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 23.485 70.035 23.555 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 14.525 70.035 14.595 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 6.685 70.035 6.755 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 291.165 70.035 291.235 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 283.325 70.035 283.395 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 275.485 70.035 275.555 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 267.645 70.035 267.715 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 259.805 70.035 259.875 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 251.965 70.035 252.035 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 244.125 70.035 244.195 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 235.165 70.035 235.235 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 228.445 70.035 228.515 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 220.605 70.035 220.675 ;
        END
    END p199
    OBS
      LAYER via2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER via1 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal1 ;
        RECT  0 0 71.54 299.04 ;
    END
END fake_macro_adaptec1_o211426

MACRO fake_macro_adaptec1_o211427
    CLASS BLOCK ;
    SIZE 71.4 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 291.165 70.035 291.235 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 283.325 70.035 283.395 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 275.485 70.035 275.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 267.645 70.035 267.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 259.805 70.035 259.875 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 251.965 70.035 252.035 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 244.125 70.035 244.195 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 235.165 70.035 235.235 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 228.445 70.035 228.515 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 220.605 70.035 220.675 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 211.645 70.035 211.715 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 204.925 70.035 204.995 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 197.085 70.035 197.155 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 188.125 70.035 188.195 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 181.405 70.035 181.475 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 173.565 70.035 173.635 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 164.605 70.035 164.675 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 157.885 70.035 157.955 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.965 70.035 140.035 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 132.125 70.035 132.195 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 124.285 70.035 124.355 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 116.445 70.035 116.515 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 108.605 70.035 108.675 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 100.765 70.035 100.835 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 94.045 70.035 94.115 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 85.085 70.035 85.155 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 77.245 70.035 77.315 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 70.525 70.035 70.595 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 61.565 70.035 61.635 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 53.725 70.035 53.795 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 47.005 70.035 47.075 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 38.045 70.035 38.115 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 30.205 70.035 30.275 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 23.485 70.035 23.555 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 14.525 70.035 14.595 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 6.685 70.035 6.755 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 153.965 68.915 154.035 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.125 69.475 153.195 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.165 0.595 144.235 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.205 68.915 142.275 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.365 3.955 148.435 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.245 2.275 147.315 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p73
    PIN p74
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p75
    PIN p76
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p77
    PIN p78
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p79
    PIN p80
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p81
    PIN p82
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p83
    PIN p84
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p85
    PIN p86
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.605 1.155 3.675 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.445 1.155 11.515 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.285 1.155 19.355 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.125 1.155 27.195 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.965 1.155 35.035 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.805 1.155 42.875 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.645 1.155 50.715 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.485 1.155 58.555 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.325 1.155 66.395 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.165 1.155 74.235 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.005 1.155 82.075 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.845 1.155 89.915 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.525 1.155 105.595 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.365 1.155 113.435 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.205 1.155 121.275 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.045 1.155 129.115 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.485 1.155 184.555 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.165 1.155 200.235 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.525 1.155 231.595 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.245 2.275 119.315 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.405 2.275 111.475 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.565 2.275 103.635 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 95.725 2.275 95.795 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 87.885 2.275 87.955 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.045 2.275 80.115 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.205 2.275 72.275 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.365 2.275 64.435 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.685 2.275 195.755 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 187.845 2.275 187.915 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.005 2.275 180.075 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.165 2.275 172.235 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.325 2.275 164.395 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.485 2.275 156.555 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.925 2.275 134.995 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.085 2.275 127.155 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.405 2.275 258.475 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.565 2.275 250.635 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 242.725 2.275 242.795 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 234.885 2.275 234.955 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.045 2.275 227.115 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.205 2.275 219.275 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.365 2.275 211.435 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.525 2.275 203.595 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 289.765 2.275 289.835 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 281.925 2.275 281.995 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.085 2.275 274.155 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.245 2.275 266.315 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 150.605 2.275 150.675 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 149.485 3.395 149.555 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.085 69.475 148.155 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.005 69.475 152.075 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 181.685 68.915 181.755 ;
        END
    END p199
    OBS
      LAYER via2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER via1 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal1 ;
        RECT  0 0 71.54 299.04 ;
    END
END fake_macro_adaptec1_o211427

MACRO fake_macro_adaptec1_o211428
    CLASS BLOCK ;
    SIZE 71.4 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 153.965 68.915 154.035 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 220.605 70.035 220.675 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 211.645 70.035 211.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 204.925 70.035 204.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 197.085 70.035 197.155 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 188.125 70.035 188.195 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 181.405 70.035 181.475 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 132.125 70.035 132.195 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 124.285 70.035 124.355 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 108.605 70.035 108.675 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 100.765 70.035 100.835 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 94.045 70.035 94.115 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 85.085 70.035 85.155 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 77.245 70.035 77.315 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 70.525 70.035 70.595 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 61.565 70.035 61.635 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 53.725 70.035 53.795 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 47.005 70.035 47.075 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 38.045 70.035 38.115 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 30.205 70.035 30.275 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 23.485 70.035 23.555 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 14.525 70.035 14.595 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 6.685 70.035 6.755 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 267.645 70.035 267.715 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 275.485 70.035 275.555 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 283.325 70.035 283.395 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 291.165 70.035 291.235 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 235.165 70.035 235.235 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 244.125 70.035 244.195 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 251.965 70.035 252.035 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 259.805 70.035 259.875 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 150.605 2.275 150.675 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.125 69.475 153.195 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.205 68.915 142.275 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.365 3.955 148.435 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.245 2.275 147.315 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 234.885 2.275 234.955 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 242.725 2.275 242.795 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.565 2.275 250.635 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.405 2.275 258.475 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.245 2.275 266.315 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 149.485 3.395 149.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.005 69.475 152.075 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 181.685 68.915 181.755 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.165 0.595 144.235 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p68
    PIN p69
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p74
    PIN p75
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.605 1.155 3.675 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.445 1.155 11.515 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.285 1.155 19.355 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.125 1.155 27.195 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.965 1.155 35.035 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.805 1.155 42.875 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.645 1.155 50.715 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.485 1.155 58.555 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.325 1.155 66.395 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.165 1.155 74.235 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.005 1.155 82.075 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.845 1.155 89.915 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.525 1.155 105.595 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.365 1.155 113.435 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.205 1.155 121.275 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.045 1.155 129.115 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.485 1.155 184.555 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.165 1.155 200.235 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.525 1.155 231.595 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.085 2.275 274.155 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 87.885 2.275 87.955 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.045 2.275 80.115 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.205 2.275 72.275 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.365 2.275 64.435 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 281.925 2.275 281.995 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.325 2.275 164.395 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.485 2.275 156.555 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.925 2.275 134.995 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.085 2.275 127.155 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.245 2.275 119.315 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.405 2.275 111.475 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.565 2.275 103.635 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 95.725 2.275 95.795 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 289.765 2.275 289.835 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.045 2.275 227.115 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.205 2.275 219.275 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.365 2.275 211.435 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.525 2.275 203.595 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.685 2.275 195.755 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 187.845 2.275 187.915 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.005 2.275 180.075 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.165 2.275 172.235 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.085 69.475 148.155 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 228.445 70.035 228.515 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 173.565 70.035 173.635 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 164.605 70.035 164.675 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 157.885 70.035 157.955 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.965 70.035 140.035 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 116.445 70.035 116.515 ;
        END
    END p199
    OBS
      LAYER via2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER via1 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal1 ;
        RECT  0 0 71.54 299.04 ;
    END
END fake_macro_adaptec1_o211428

MACRO fake_macro_adaptec1_o211429
    CLASS BLOCK ;
    SIZE 71.4 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 291.165 70.035 291.235 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 283.325 70.035 283.395 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 275.485 70.035 275.555 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 267.645 70.035 267.715 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 259.805 70.035 259.875 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 251.965 70.035 252.035 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 235.165 70.035 235.235 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 228.445 70.035 228.515 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 220.605 70.035 220.675 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 211.645 70.035 211.715 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 204.925 70.035 204.995 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 197.085 70.035 197.155 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 188.125 70.035 188.195 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 181.405 70.035 181.475 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 173.565 70.035 173.635 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 164.605 70.035 164.675 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 157.885 70.035 157.955 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.965 70.035 140.035 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 132.125 70.035 132.195 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 124.285 70.035 124.355 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 116.445 70.035 116.515 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 108.605 70.035 108.675 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 100.765 70.035 100.835 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 94.045 70.035 94.115 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 85.085 70.035 85.155 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 77.245 70.035 77.315 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 70.525 70.035 70.595 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 61.565 70.035 61.635 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 53.725 70.035 53.795 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 47.005 70.035 47.075 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 38.045 70.035 38.115 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 30.205 70.035 30.275 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 23.485 70.035 23.555 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 14.525 70.035 14.595 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 6.685 70.035 6.755 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 153.965 68.915 154.035 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.125 69.475 153.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.205 68.915 142.275 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.365 3.955 148.435 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.245 2.275 147.315 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 150.605 2.275 150.675 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 149.485 3.395 149.555 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.085 69.475 148.155 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.005 69.475 152.075 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 181.685 68.915 181.755 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.165 0.595 144.235 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p68
    PIN p69
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p74
    PIN p75
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.605 1.155 3.675 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.445 1.155 11.515 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.285 1.155 19.355 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.125 1.155 27.195 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.965 1.155 35.035 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.805 1.155 42.875 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.645 1.155 50.715 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.485 1.155 58.555 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.325 1.155 66.395 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.165 1.155 74.235 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.005 1.155 82.075 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.845 1.155 89.915 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.525 1.155 105.595 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.365 1.155 113.435 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.205 1.155 121.275 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.045 1.155 129.115 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.485 1.155 184.555 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.165 1.155 200.235 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.525 1.155 231.595 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.245 2.275 119.315 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.405 2.275 111.475 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.565 2.275 103.635 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 95.725 2.275 95.795 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 87.885 2.275 87.955 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.045 2.275 80.115 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.205 2.275 72.275 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.365 2.275 64.435 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.685 2.275 195.755 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 187.845 2.275 187.915 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.005 2.275 180.075 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.165 2.275 172.235 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.325 2.275 164.395 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.485 2.275 156.555 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.925 2.275 134.995 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.085 2.275 127.155 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.405 2.275 258.475 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.565 2.275 250.635 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 242.725 2.275 242.795 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 234.885 2.275 234.955 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.045 2.275 227.115 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.205 2.275 219.275 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.365 2.275 211.435 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.525 2.275 203.595 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 289.765 2.275 289.835 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 281.925 2.275 281.995 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.085 2.275 274.155 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.245 2.275 266.315 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 244.125 70.035 244.195 ;
        END
    END p199
    OBS
      LAYER via2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER via1 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal1 ;
        RECT  0 0 71.54 299.04 ;
    END
END fake_macro_adaptec1_o211429

MACRO fake_macro_adaptec1_o211430
    CLASS BLOCK ;
    SIZE 71.4 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p0
    PIN p1
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 228.445 70.035 228.515 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 220.605 70.035 220.675 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 211.645 70.035 211.715 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 204.925 70.035 204.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 197.085 70.035 197.155 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 181.405 70.035 181.475 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 173.565 70.035 173.635 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 164.605 70.035 164.675 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 157.885 70.035 157.955 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 139.965 70.035 140.035 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 132.125 70.035 132.195 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 124.285 70.035 124.355 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 116.445 70.035 116.515 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 108.605 70.035 108.675 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 100.765 70.035 100.835 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 94.045 70.035 94.115 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 85.085 70.035 85.155 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 77.245 70.035 77.315 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 70.525 70.035 70.595 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 61.565 70.035 61.635 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 53.725 70.035 53.795 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 47.005 70.035 47.075 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 38.045 70.035 38.115 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 30.205 70.035 30.275 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 23.485 70.035 23.555 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 14.525 70.035 14.595 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 6.685 70.035 6.755 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 267.645 70.035 267.715 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 275.485 70.035 275.555 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 283.325 70.035 283.395 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 291.165 70.035 291.235 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 235.165 70.035 235.235 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 244.125 70.035 244.195 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 251.965 70.035 252.035 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 259.805 70.035 259.875 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 150.605 2.275 150.675 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 153.965 68.915 154.035 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 153.125 69.475 153.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 142.485 69.475 142.555 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 142.205 68.915 142.275 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.885 148.365 3.955 148.435 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 147.245 2.275 147.315 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  3.325 149.485 3.395 149.555 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 148.085 69.475 148.155 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 152.005 69.475 152.075 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.765 0.595 142.835 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 144.165 0.595 144.235 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 234.885 2.275 234.955 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 242.725 2.275 242.795 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 250.565 2.275 250.635 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 258.405 2.275 258.475 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 266.245 2.275 266.315 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 239.365 1.155 239.435 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 247.205 1.155 247.275 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 255.045 1.155 255.115 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 262.885 1.155 262.955 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 270.725 1.155 270.795 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 278.565 1.155 278.635 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 286.405 1.155 286.475 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 294.245 1.155 294.315 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 3.605 1.155 3.675 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 11.445 1.155 11.515 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 19.285 1.155 19.355 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 27.125 1.155 27.195 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 34.965 1.155 35.035 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 42.805 1.155 42.875 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 50.645 1.155 50.715 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 58.485 1.155 58.555 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.325 1.155 66.395 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 74.165 1.155 74.235 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 82.005 1.155 82.075 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 89.845 1.155 89.915 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 97.685 1.155 97.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 105.525 1.155 105.595 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 113.365 1.155 113.435 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 121.205 1.155 121.275 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 129.045 1.155 129.115 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 136.885 1.155 136.955 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 160.965 1.155 161.035 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 168.805 1.155 168.875 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 176.645 1.155 176.715 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 184.485 1.155 184.555 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 192.325 1.155 192.395 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 200.165 1.155 200.235 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 208.005 1.155 208.075 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 215.845 1.155 215.915 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 223.685 1.155 223.755 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 231.525 1.155 231.595 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 274.085 2.275 274.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 87.885 2.275 87.955 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 80.045 2.275 80.115 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 72.205 2.275 72.275 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 64.365 2.275 64.435 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 164.325 2.275 164.395 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 156.485 2.275 156.555 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 134.925 2.275 134.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 127.085 2.275 127.155 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 119.245 2.275 119.315 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 111.405 2.275 111.475 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 103.565 2.275 103.635 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 95.725 2.275 95.795 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 172.165 2.275 172.235 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 289.765 2.275 289.835 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 227.045 2.275 227.115 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 219.205 2.275 219.275 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 211.365 2.275 211.435 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 203.525 2.275 203.595 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 195.685 2.275 195.755 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 187.845 2.275 187.915 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 180.005 2.275 180.075 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 281.925 2.275 281.995 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 172.725 0.595 172.795 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.085 0.595 204.155 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 258.965 0.595 259.035 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 181.685 68.915 181.755 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 188.125 70.035 188.195 ;
        END
    END p199
    OBS
      LAYER via2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal2 ;
        RECT  0 0 71.54 299.04 ;
      LAYER via1 ;
        RECT  0 0 71.54 299.04 ;
      LAYER metal1 ;
        RECT  0 0 71.54 299.04 ;
    END
END fake_macro_adaptec1_o211430

MACRO fake_macro_adaptec1_o211431
    CLASS BLOCK ;
    SIZE 38.64 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 152.005 36.995 152.075 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 153.965 36.995 154.035 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 181.685 36.995 181.755 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 153.685 36.995 153.755 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 142.205 36.995 142.275 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 153.405 36.995 153.475 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 9.765 0.595 9.835 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 56.805 0.595 56.875 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.325 0.595 192.395 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 168.805 0.595 168.875 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 262.885 0.595 262.955 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.365 0.595 239.435 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 215.845 0.595 215.915 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.245 0.595 294.315 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.405 0.595 286.475 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p87
    PIN p88
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 53.725 36.995 53.795 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 49.805 36.995 49.875 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 45.885 36.995 45.955 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 41.965 36.995 42.035 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 38.045 36.995 38.115 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 34.125 36.995 34.195 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 30.205 36.995 30.275 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 26.285 36.995 26.355 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 22.365 36.995 22.435 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 18.445 36.995 18.515 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 14.525 36.995 14.595 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 10.605 36.995 10.675 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 6.685 36.995 6.755 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 2.765 36.995 2.835 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 295.085 36.995 295.155 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 291.165 36.995 291.235 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 287.245 36.995 287.315 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 283.325 36.995 283.395 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 279.405 36.995 279.475 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 275.485 36.995 275.555 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 271.565 36.995 271.635 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 267.645 36.995 267.715 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 263.725 36.995 263.795 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 259.805 36.995 259.875 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 255.885 36.995 255.955 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 251.965 36.995 252.035 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 224.525 36.995 224.595 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 248.045 36.995 248.115 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 220.605 36.995 220.675 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 244.125 36.995 244.195 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 216.685 36.995 216.755 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 240.205 36.995 240.275 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 212.765 36.995 212.835 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 236.285 36.995 236.355 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 208.845 36.995 208.915 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 232.365 36.995 232.435 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 204.925 36.995 204.995 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 228.445 36.995 228.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 201.005 36.995 201.075 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 197.085 36.995 197.155 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 193.165 36.995 193.235 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 189.245 36.995 189.315 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 185.325 36.995 185.395 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 181.405 36.995 181.475 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 177.485 36.995 177.555 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 173.565 36.995 173.635 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 169.645 36.995 169.715 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 165.725 36.995 165.795 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 161.805 36.995 161.875 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 157.885 36.995 157.955 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 139.965 36.995 140.035 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 136.045 36.995 136.115 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 132.125 36.995 132.195 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 128.205 36.995 128.275 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 124.285 36.995 124.355 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 120.365 36.995 120.435 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 116.445 36.995 116.515 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 112.525 36.995 112.595 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 108.605 36.995 108.675 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 104.685 36.995 104.755 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 100.765 36.995 100.835 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 96.845 36.995 96.915 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 92.925 36.995 92.995 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 89.005 36.995 89.075 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 85.085 36.995 85.155 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 81.165 36.995 81.235 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 77.245 36.995 77.315 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 73.325 36.995 73.395 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 69.405 36.995 69.475 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 65.485 36.995 65.555 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 61.565 36.995 61.635 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 57.645 36.995 57.715 ;
        END
    END p375
    OBS
      LAYER via2 ;
        RECT  0 0 38.64 299.04 ;
      LAYER metal2 ;
        RECT  0 0 38.64 299.04 ;
      LAYER via1 ;
        RECT  0 0 38.64 299.04 ;
      LAYER metal1 ;
        RECT  0 0 38.64 299.04 ;
    END
END fake_macro_adaptec1_o211431

MACRO fake_macro_adaptec1_o211432
    CLASS BLOCK ;
    SIZE 38.64 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 149.485 1.715 149.555 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 152.005 36.995 152.075 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 153.965 36.995 154.035 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 181.685 36.995 181.755 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 153.685 36.995 153.755 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 142.205 36.995 142.275 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 153.405 36.995 153.475 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.645 148.365 1.715 148.435 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 148.365 2.835 148.435 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.765 149.485 2.835 149.555 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.565 0.595 68.635 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 56.805 0.595 56.875 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.125 0.595 41.195 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.685 0.595 13.755 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 9.765 0.595 9.835 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.165 0.595 200.235 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.325 0.595 192.395 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.565 0.595 180.635 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 168.805 0.595 168.875 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.365 0.595 239.435 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.605 0.595 227.675 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 215.845 0.595 215.915 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.005 0.595 208.075 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.245 0.595 294.315 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.405 0.595 286.475 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.485 0.595 282.555 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.645 0.595 274.715 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 262.885 0.595 262.955 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.045 0.595 255.115 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.885 0.595 248.955 ;
        END
    END p89
    PIN p90
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 14.525 36.995 14.595 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 10.605 36.995 10.675 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 6.685 36.995 6.755 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 2.765 36.995 2.835 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 287.245 36.995 287.315 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 283.325 36.995 283.395 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 279.405 36.995 279.475 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 275.485 36.995 275.555 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 271.565 36.995 271.635 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 267.645 36.995 267.715 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 224.525 36.995 224.595 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 220.605 36.995 220.675 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 216.685 36.995 216.755 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 212.765 36.995 212.835 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 208.845 36.995 208.915 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 204.925 36.995 204.995 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 201.005 36.995 201.075 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 197.085 36.995 197.155 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 193.165 36.995 193.235 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 189.245 36.995 189.315 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 185.325 36.995 185.395 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 181.405 36.995 181.475 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 177.485 36.995 177.555 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 173.565 36.995 173.635 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 169.645 36.995 169.715 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 165.725 36.995 165.795 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 161.805 36.995 161.875 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 157.885 36.995 157.955 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 139.965 36.995 140.035 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 136.045 36.995 136.115 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 132.125 36.995 132.195 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 128.205 36.995 128.275 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 124.285 36.995 124.355 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 120.365 36.995 120.435 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 116.445 36.995 116.515 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 112.525 36.995 112.595 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 108.605 36.995 108.675 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 104.685 36.995 104.755 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 100.765 36.995 100.835 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 96.845 36.995 96.915 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 92.925 36.995 92.995 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 89.005 36.995 89.075 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 85.085 36.995 85.155 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 81.165 36.995 81.235 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 77.245 36.995 77.315 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 73.325 36.995 73.395 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 69.405 36.995 69.475 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 65.485 36.995 65.555 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 61.565 36.995 61.635 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 57.645 36.995 57.715 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 295.085 36.995 295.155 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 291.165 36.995 291.235 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 263.725 36.995 263.795 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 259.805 36.995 259.875 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 255.885 36.995 255.955 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 251.965 36.995 252.035 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 248.045 36.995 248.115 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 244.125 36.995 244.195 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 240.205 36.995 240.275 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 236.285 36.995 236.355 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 232.365 36.995 232.435 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 228.445 36.995 228.515 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 53.725 36.995 53.795 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 49.805 36.995 49.875 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 45.885 36.995 45.955 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 41.965 36.995 42.035 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 38.045 36.995 38.115 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 34.125 36.995 34.195 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 30.205 36.995 30.275 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 26.285 36.995 26.355 ;
        END
    END p373
    PIN p374
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 22.365 36.995 22.435 ;
        END
    END p374
    PIN p375
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  36.925 18.445 36.995 18.515 ;
        END
    END p375
    OBS
      LAYER via2 ;
        RECT  0 0 38.64 299.04 ;
      LAYER metal2 ;
        RECT  0 0 38.64 299.04 ;
      LAYER via1 ;
        RECT  0 0 38.64 299.04 ;
      LAYER metal1 ;
        RECT  0 0 38.64 299.04 ;
    END
END fake_macro_adaptec1_o211432

MACRO fake_macro_adaptec1_o211433
    CLASS BLOCK ;
    SIZE 11.2 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.245 0.595 294.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.405 0.595 286.475 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 262.885 0.595 262.955 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.805 0.595 252.875 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.365 0.595 239.435 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.205 0.595 233.275 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 215.845 0.595 215.915 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.325 0.595 192.395 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.325 0.595 178.395 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 168.805 0.595 168.875 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.725 0.595 158.795 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.085 0.595 141.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.485 0.595 121.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 56.805 0.595 56.875 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 9.765 0.595 9.835 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 152.005 9.555 152.075 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 142.205 9.555 142.275 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 169.925 9.555 169.995 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 153.965 9.555 154.035 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 153.685 9.555 153.755 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 85.085 9.555 85.155 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 81.165 9.555 81.235 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 77.245 9.555 77.315 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 73.325 9.555 73.395 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 69.405 9.555 69.475 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 65.485 9.555 65.555 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 61.565 9.555 61.635 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 57.645 9.555 57.715 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 53.725 9.555 53.795 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 49.805 9.555 49.875 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 45.885 9.555 45.955 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 38.045 9.555 38.115 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 34.125 9.555 34.195 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 30.205 9.555 30.275 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 26.285 9.555 26.355 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 22.365 9.555 22.435 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 18.445 9.555 18.515 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 14.525 9.555 14.595 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.605 9.555 10.675 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 6.685 9.555 6.755 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.765 9.555 2.835 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 255.885 9.555 255.955 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 251.965 9.555 252.035 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 248.045 9.555 248.115 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 244.125 9.555 244.195 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 240.205 9.555 240.275 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 236.285 9.555 236.355 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 232.365 9.555 232.435 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 228.445 9.555 228.515 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 224.525 9.555 224.595 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 220.605 9.555 220.675 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 216.685 9.555 216.755 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 212.765 9.555 212.835 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 208.845 9.555 208.915 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 204.925 9.555 204.995 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 201.005 9.555 201.075 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 197.085 9.555 197.155 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 193.165 9.555 193.235 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 189.245 9.555 189.315 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 185.325 9.555 185.395 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 181.405 9.555 181.475 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 295.085 9.555 295.155 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 291.165 9.555 291.235 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 287.245 9.555 287.315 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 283.325 9.555 283.395 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 279.405 9.555 279.475 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 275.485 9.555 275.555 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 271.565 9.555 271.635 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 177.485 9.555 177.555 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 267.645 9.555 267.715 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 173.565 9.555 173.635 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 263.725 9.555 263.795 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 169.645 9.555 169.715 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 259.805 9.555 259.875 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 165.725 9.555 165.795 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 161.805 9.555 161.875 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 157.885 9.555 157.955 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 139.965 9.555 140.035 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 136.045 9.555 136.115 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 132.125 9.555 132.195 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.205 9.555 128.275 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 124.285 9.555 124.355 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 120.365 9.555 120.435 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 116.445 9.555 116.515 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 112.525 9.555 112.595 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 108.605 9.555 108.675 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 104.685 9.555 104.755 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 100.765 9.555 100.835 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 96.845 9.555 96.915 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 92.925 9.555 92.995 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 89.005 9.555 89.075 ;
        END
    END p369
    OBS
      LAYER via2 ;
        RECT  0 0 11.2 299.04 ;
      LAYER metal2 ;
        RECT  0 0 11.2 299.04 ;
      LAYER via1 ;
        RECT  0 0 11.2 299.04 ;
      LAYER metal1 ;
        RECT  0 0 11.2 299.04 ;
    END
END fake_macro_adaptec1_o211433

MACRO fake_macro_adaptec1_o211434
    CLASS BLOCK ;
    SIZE 11.2 BY 142.8 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 75.565 9.555 75.635 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.445 0.595 123.515 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.845 0.595 117.915 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.605 0.595 115.675 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.005 0.595 110.075 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.085 0.595 106.155 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.005 0.595 96.075 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.085 0.595 92.155 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.165 0.595 88.235 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.565 0.595 82.635 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.685 0.595 62.755 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 56.805 0.595 56.875 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.405 0.595 27.475 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.525 0.595 21.595 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 103.285 9.555 103.355 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 137.725 0.595 137.795 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 73.605 9.555 73.675 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 75.285 9.555 75.355 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p68
    PIN p69
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.045 0.595 80.115 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.965 0.595 84.035 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.925 0.595 78.995 ;
        END
    END p74
    PIN p75
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.885 0.595 87.955 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.845 0.595 82.915 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.805 0.595 91.875 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.765 0.595 86.835 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.725 0.595 95.795 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.685 0.595 90.755 ;
        END
    END p80
    PIN p81
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.645 0.595 99.715 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.605 0.595 94.675 ;
        END
    END p82
    PIN p83
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.565 0.595 103.635 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 98.525 0.595 98.595 ;
        END
    END p84
    PIN p85
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.485 0.595 107.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 102.445 0.595 102.515 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.405 0.595 111.475 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.365 0.595 106.435 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.325 0.595 115.395 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.285 0.595 110.355 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.245 0.595 119.315 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.205 0.595 114.275 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.165 0.595 123.235 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.125 0.595 118.195 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.085 0.595 127.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.045 0.595 122.115 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.005 0.595 131.075 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.965 0.595 126.035 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.925 0.595 134.995 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.885 0.595 129.955 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.845 0.595 138.915 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.805 0.595 133.875 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 79.485 0.595 79.555 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.405 0.595 83.475 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.325 0.595 87.395 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.245 0.595 91.315 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.165 0.595 95.235 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.085 0.595 99.155 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.005 0.595 103.075 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 106.925 0.595 106.995 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 110.845 0.595 110.915 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 114.765 0.595 114.835 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.685 0.595 118.755 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.605 0.595 122.675 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.525 0.595 126.595 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.445 0.595 130.515 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.365 0.595 134.435 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.285 0.595 138.355 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 63.805 9.555 63.875 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 75.005 9.555 75.075 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 99.085 9.555 99.155 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 95.165 9.555 95.235 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 91.245 9.555 91.315 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 87.325 9.555 87.395 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 83.405 9.555 83.475 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 79.485 9.555 79.555 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 61.565 9.555 61.635 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 57.645 9.555 57.715 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 53.725 9.555 53.795 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 49.805 9.555 49.875 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 45.885 9.555 45.955 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 38.045 9.555 38.115 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 34.125 9.555 34.195 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 30.205 9.555 30.275 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 26.285 9.555 26.355 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 22.365 9.555 22.435 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 18.445 9.555 18.515 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 14.525 9.555 14.595 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.605 9.555 10.675 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 6.685 9.555 6.755 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.765 9.555 2.835 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 138.285 9.555 138.355 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 134.365 9.555 134.435 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 130.445 9.555 130.515 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 126.525 9.555 126.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 122.605 9.555 122.675 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 118.685 9.555 118.755 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 114.765 9.555 114.835 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 110.845 9.555 110.915 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 106.925 9.555 106.995 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 103.005 9.555 103.075 ;
        END
    END p169
    OBS
      LAYER via2 ;
        RECT  0 0 11.2 142.8 ;
      LAYER metal2 ;
        RECT  0 0 11.2 142.8 ;
      LAYER via1 ;
        RECT  0 0 11.2 142.8 ;
      LAYER metal1 ;
        RECT  0 0 11.2 142.8 ;
    END
END fake_macro_adaptec1_o211434

MACRO fake_macro_adaptec1_o211435
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.685 21.315 181.755 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.405 21.315 153.475 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p303
    PIN p304
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p304
    PIN p305
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p305
    PIN p306
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p306
    PIN p307
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p307
    PIN p308
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p308
    PIN p309
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p309
    PIN p310
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p310
    PIN p311
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p311
    PIN p312
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p312
    PIN p313
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p313
    PIN p314
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p314
    PIN p315
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p315
    PIN p316
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p316
    PIN p317
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p317
    PIN p318
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p318
    PIN p319
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p319
    PIN p320
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p320
    PIN p321
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p321
    PIN p322
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p322
    PIN p323
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p323
    PIN p324
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p324
    PIN p325
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p325
    PIN p326
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p326
    PIN p327
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p327
    PIN p328
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p329
    PIN p330
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o211435

MACRO fake_macro_adaptec1_o211436
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p1
    PIN p2
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.685 21.315 181.755 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.405 21.315 153.475 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p303
    PIN p304
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p304
    PIN p305
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p305
    PIN p306
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p306
    PIN p307
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p307
    PIN p308
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p308
    PIN p309
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p309
    PIN p310
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p310
    PIN p311
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p311
    PIN p312
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p312
    PIN p313
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p313
    PIN p314
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p314
    PIN p315
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p315
    PIN p316
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p316
    PIN p317
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p317
    PIN p318
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p318
    PIN p319
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p319
    PIN p320
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p320
    PIN p321
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p321
    PIN p322
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p322
    PIN p323
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p323
    PIN p324
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p324
    PIN p325
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p325
    PIN p326
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p326
    PIN p327
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p327
    PIN p328
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p329
    PIN p330
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o211436

MACRO fake_macro_adaptec1_o211437
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.925 21.315 169.995 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 154.245 21.875 154.315 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p88
    PIN p89
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p90
    PIN p91
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o211437

MACRO fake_macro_adaptec1_o211438
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p68
    PIN p69
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p73
    PIN p74
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p74
    PIN p75
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p78
    PIN p79
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.685 21.315 181.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.405 21.315 153.475 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p123
    PIN p124
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p125
    PIN p126
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p127
    PIN p128
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p129
    PIN p130
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p131
    PIN p132
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p133
    PIN p134
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p135
    PIN p136
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p137
    PIN p138
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p139
    PIN p140
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p141
    PIN p142
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p143
    PIN p144
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p145
    PIN p146
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p147
    PIN p148
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p149
    PIN p150
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p151
    PIN p152
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p153
    PIN p154
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p155
    PIN p156
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p157
    PIN p158
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p303
    PIN p304
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p304
    PIN p305
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p305
    PIN p306
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p306
    PIN p307
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p307
    PIN p308
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p308
    PIN p309
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p309
    PIN p310
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p310
    PIN p311
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p311
    PIN p312
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p312
    PIN p313
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p313
    PIN p314
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p314
    PIN p315
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p315
    PIN p316
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p316
    PIN p317
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p317
    PIN p318
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p318
    PIN p319
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p319
    PIN p320
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p320
    PIN p321
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p321
    PIN p322
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p322
    PIN p323
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p323
    PIN p324
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p324
    PIN p325
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p325
    PIN p326
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p326
    PIN p327
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p327
    PIN p328
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p329
    PIN p330
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p330
    PIN p331
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p331
    PIN p332
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p332
    PIN p333
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p333
    PIN p334
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p334
    PIN p335
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p335
    PIN p336
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p336
    PIN p337
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p337
    PIN p338
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p338
    PIN p339
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p339
    PIN p340
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p340
    PIN p341
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p341
    PIN p342
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p342
    PIN p343
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p343
    PIN p344
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p344
    PIN p345
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p345
    PIN p346
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p346
    PIN p347
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p347
    PIN p348
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p348
    PIN p349
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p349
    PIN p350
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p350
    PIN p351
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p351
    PIN p352
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p352
    PIN p353
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p353
    PIN p354
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p354
    PIN p355
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p355
    PIN p356
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p356
    PIN p357
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p357
    PIN p358
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p358
    PIN p359
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p359
    PIN p360
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p360
    PIN p361
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p361
    PIN p362
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p362
    PIN p363
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p363
    PIN p364
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p364
    PIN p365
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p365
    PIN p366
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p366
    PIN p367
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p367
    PIN p368
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p368
    PIN p369
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p369
    PIN p370
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p370
    PIN p371
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p371
    PIN p372
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p372
    PIN p373
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o211438

MACRO fake_macro_adaptec1_o211439
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p2
    PIN p3
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p3
    PIN p4
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p4
    PIN p5
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p5
    PIN p6
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p6
    PIN p7
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p7
    PIN p8
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p8
    PIN p9
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p9
    PIN p10
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p11
    PIN p12
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p12
    PIN p13
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p13
    PIN p14
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p14
    PIN p15
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p20
    PIN p21
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p39
    PIN p40
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p41
    PIN p42
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p43
    PIN p44
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p45
    PIN p46
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p47
    PIN p48
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p49
    PIN p50
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p50
    PIN p51
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p51
    PIN p52
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p52
    PIN p53
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p53
    PIN p54
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p54
    PIN p55
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p55
    PIN p56
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p56
    PIN p57
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p57
    PIN p58
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p58
    PIN p59
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p59
    PIN p60
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p60
    PIN p61
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p61
    PIN p62
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p62
    PIN p63
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p63
    PIN p64
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p64
    PIN p65
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p65
    PIN p66
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p66
    PIN p67
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p67
    PIN p68
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p68
    PIN p69
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p70
    PIN p71
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p71
    PIN p72
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p72
    PIN p73
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p73
    PIN p74
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p76
    PIN p77
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.925 21.315 169.995 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p124
    PIN p125
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p126
    PIN p127
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p128
    PIN p129
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p130
    PIN p131
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p132
    PIN p133
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p134
    PIN p135
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p136
    PIN p137
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p138
    PIN p139
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p140
    PIN p141
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p142
    PIN p143
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p144
    PIN p145
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p146
    PIN p147
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p148
    PIN p149
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p150
    PIN p151
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p152
    PIN p153
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p297
    PIN p298
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p299
    PIN p300
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 154.245 21.875 154.315 ;
        END
    END p301
    PIN p302
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p302
    PIN p303
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p303
    PIN p304
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p304
    PIN p305
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p305
    PIN p306
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p306
    PIN p307
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p307
    PIN p308
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p308
    PIN p309
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p309
    PIN p310
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p310
    PIN p311
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p311
    PIN p312
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p312
    PIN p313
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p313
    PIN p314
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p314
    PIN p315
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p315
    PIN p316
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p316
    PIN p317
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p317
    PIN p318
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p318
    PIN p319
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p319
    PIN p320
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p320
    PIN p321
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p321
    PIN p322
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p322
    PIN p323
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p323
    PIN p324
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p324
    PIN p325
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p325
    PIN p326
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p326
    PIN p327
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p327
    PIN p328
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p328
    PIN p329
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p329
    PIN p330
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p330
    PIN p331
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p331
    PIN p332
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p332
    PIN p333
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p333
    PIN p334
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p334
    PIN p335
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p335
    PIN p336
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p336
    PIN p337
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p337
    PIN p338
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p338
    PIN p339
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p339
    PIN p340
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p340
    PIN p341
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p341
    PIN p342
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p342
    PIN p343
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p343
    PIN p344
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p344
    PIN p345
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p345
    PIN p346
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p346
    PIN p347
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p347
    PIN p348
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p348
    PIN p349
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p349
    PIN p350
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p350
    PIN p351
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p351
    PIN p352
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p352
    PIN p353
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p353
    PIN p354
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p354
    PIN p355
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p355
    PIN p356
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p356
    PIN p357
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p357
    PIN p358
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p358
    PIN p359
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p359
    PIN p360
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p360
    PIN p361
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p361
    PIN p362
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p362
    PIN p363
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p363
    PIN p364
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p364
    PIN p365
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p365
    PIN p366
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p366
    PIN p367
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p367
    PIN p368
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p368
    PIN p369
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p369
    PIN p370
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p370
    PIN p371
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p371
    PIN p372
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p372
    PIN p373
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o211439

MACRO fake_macro_adaptec1_o211440
    CLASS BLOCK ;
    SIZE 22.96 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 142.205 21.315 142.275 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.925 21.315 169.995 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.965 21.315 154.035 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 148.365 2.275 148.435 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 148.365 0.595 148.435 ;
        END
    END p69
    PIN p70
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.805 154.245 21.875 154.315 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 153.685 21.315 153.755 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 152.005 21.315 152.075 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 149.485 0.595 149.555 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 149.485 2.275 149.555 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.485 0.595 268.555 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.325 0.595 31.395 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.725 0.595 11.795 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.805 0.595 7.875 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.885 0.595 3.955 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.765 0.595 58.835 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.845 0.595 54.915 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.045 0.595 45.115 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 35.245 0.595 35.315 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 86.205 0.595 86.275 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.285 0.595 82.355 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.645 0.595 64.715 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.525 0.595 119.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.725 0.595 109.795 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.805 0.595 105.875 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.885 0.595 101.955 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.485 0.595 170.555 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.565 0.595 166.635 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.045 0.595 157.115 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.125 0.595 139.195 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 133.245 0.595 133.315 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.325 0.595 129.395 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 288.085 0.595 288.155 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.925 0.595 197.995 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 194.005 0.595 194.075 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 190.085 0.595 190.155 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.645 0.595 176.715 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 292.005 0.595 292.075 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.525 0.595 231.595 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.445 0.595 221.515 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.525 0.595 217.595 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.605 0.595 213.675 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.925 0.595 295.995 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.565 0.595 264.635 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p154
    PIN p155
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.125 0.595 251.195 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p156
    PIN p157
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.965 0.595 245.035 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 241.045 0.595 241.115 ;
        END
    END p158
    PIN p159
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p159
    PIN p160
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p160
    PIN p161
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p161
    PIN p162
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p162
    PIN p163
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p163
    PIN p164
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p164
    PIN p165
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p165
    PIN p166
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p166
    PIN p167
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p167
    PIN p168
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p168
    PIN p169
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p169
    PIN p170
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p170
    PIN p171
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p171
    PIN p172
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p172
    PIN p173
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p173
    PIN p174
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p174
    PIN p175
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p175
    PIN p176
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p176
    PIN p177
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p177
    PIN p178
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p178
    PIN p179
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p179
    PIN p180
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p180
    PIN p181
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p181
    PIN p182
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p182
    PIN p183
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p183
    PIN p184
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p184
    PIN p185
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p185
    PIN p186
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p186
    PIN p187
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p187
    PIN p188
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p188
    PIN p189
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p189
    PIN p190
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p190
    PIN p191
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p191
    PIN p192
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p192
    PIN p193
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p193
    PIN p194
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p194
    PIN p195
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p195
    PIN p196
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p196
    PIN p197
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p197
    PIN p198
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p198
    PIN p199
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p199
    PIN p200
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p200
    PIN p201
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p201
    PIN p202
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p202
    PIN p203
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p203
    PIN p204
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p204
    PIN p205
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p205
    PIN p206
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p206
    PIN p207
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p207
    PIN p208
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p208
    PIN p209
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p209
    PIN p210
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p210
    PIN p211
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p211
    PIN p212
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p212
    PIN p213
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p213
    PIN p214
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p214
    PIN p215
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p215
    PIN p216
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p216
    PIN p217
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p217
    PIN p218
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p218
    PIN p219
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p219
    PIN p220
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p220
    PIN p221
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p221
    PIN p222
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p222
    PIN p223
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p223
    PIN p224
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p224
    PIN p225
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p225
    PIN p226
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p226
    PIN p227
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p227
    PIN p228
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p228
    PIN p229
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p229
    PIN p230
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p230
    PIN p231
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p231
    PIN p232
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p232
    PIN p233
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p233
    PIN p234
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p234
    PIN p235
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p235
    PIN p236
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p236
    PIN p237
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p237
    PIN p238
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p238
    PIN p239
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p239
    PIN p240
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p240
    PIN p241
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p241
    PIN p242
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p242
    PIN p243
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p243
    PIN p244
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p244
    PIN p245
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p245
    PIN p246
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p246
    PIN p247
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p247
    PIN p248
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p248
    PIN p249
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p249
    PIN p250
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p250
    PIN p251
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p251
    PIN p252
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p252
    PIN p253
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p253
    PIN p254
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p254
    PIN p255
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p255
    PIN p256
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p256
    PIN p257
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p257
    PIN p258
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p258
    PIN p259
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p259
    PIN p260
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p260
    PIN p261
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p261
    PIN p262
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p262
    PIN p263
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p263
    PIN p264
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p264
    PIN p265
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p265
    PIN p266
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p266
    PIN p267
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p267
    PIN p268
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p268
    PIN p269
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p269
    PIN p270
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p270
    PIN p271
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p271
    PIN p272
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p272
    PIN p273
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p273
    PIN p274
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p274
    PIN p275
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p275
    PIN p276
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p276
    PIN p277
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p277
    PIN p278
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p278
    PIN p279
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p279
    PIN p280
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p280
    PIN p281
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p281
    PIN p282
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p282
    PIN p283
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p283
    PIN p284
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p284
    PIN p285
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p285
    PIN p286
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p286
    PIN p287
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p287
    PIN p288
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p288
    PIN p289
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p289
    PIN p290
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p290
    PIN p291
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p291
    PIN p292
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p292
    PIN p293
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p293
    PIN p294
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p294
    PIN p295
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p295
    PIN p296
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p296
    PIN p297
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p298
    PIN p299
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p300
    PIN p301
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 85.085 21.315 85.155 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 81.165 21.315 81.235 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 77.245 21.315 77.315 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 73.325 21.315 73.395 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 69.405 21.315 69.475 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 65.485 21.315 65.555 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 61.565 21.315 61.635 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 57.645 21.315 57.715 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 53.725 21.315 53.795 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 49.805 21.315 49.875 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 45.885 21.315 45.955 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 41.965 21.315 42.035 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 38.045 21.315 38.115 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 34.125 21.315 34.195 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 30.205 21.315 30.275 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 26.285 21.315 26.355 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 22.365 21.315 22.435 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 18.445 21.315 18.515 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 14.525 21.315 14.595 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 10.605 21.315 10.675 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 6.685 21.315 6.755 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 2.765 21.315 2.835 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 255.885 21.315 255.955 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 251.965 21.315 252.035 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 248.045 21.315 248.115 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 244.125 21.315 244.195 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 240.205 21.315 240.275 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 236.285 21.315 236.355 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 232.365 21.315 232.435 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 228.445 21.315 228.515 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 224.525 21.315 224.595 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 220.605 21.315 220.675 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 216.685 21.315 216.755 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 212.765 21.315 212.835 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 208.845 21.315 208.915 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 204.925 21.315 204.995 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 201.005 21.315 201.075 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 197.085 21.315 197.155 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 193.165 21.315 193.235 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 189.245 21.315 189.315 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 185.325 21.315 185.395 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 181.405 21.315 181.475 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 177.485 21.315 177.555 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 173.565 21.315 173.635 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 169.645 21.315 169.715 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 165.725 21.315 165.795 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 161.805 21.315 161.875 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 157.885 21.315 157.955 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 139.965 21.315 140.035 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 136.045 21.315 136.115 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 132.125 21.315 132.195 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 128.205 21.315 128.275 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 124.285 21.315 124.355 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 120.365 21.315 120.435 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 116.445 21.315 116.515 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 112.525 21.315 112.595 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 108.605 21.315 108.675 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 104.685 21.315 104.755 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 100.765 21.315 100.835 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 96.845 21.315 96.915 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 92.925 21.315 92.995 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 89.005 21.315 89.075 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 295.085 21.315 295.155 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 291.165 21.315 291.235 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 287.245 21.315 287.315 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 283.325 21.315 283.395 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 279.405 21.315 279.475 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 275.485 21.315 275.555 ;
        END
    END p369
    PIN p370
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 271.565 21.315 271.635 ;
        END
    END p370
    PIN p371
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 267.645 21.315 267.715 ;
        END
    END p371
    PIN p372
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 263.725 21.315 263.795 ;
        END
    END p372
    PIN p373
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  21.245 259.805 21.315 259.875 ;
        END
    END p373
    OBS
      LAYER via2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal2 ;
        RECT  0 0 22.96 299.04 ;
      LAYER via1 ;
        RECT  0 0 22.96 299.04 ;
      LAYER metal1 ;
        RECT  0 0 22.96 299.04 ;
    END
END fake_macro_adaptec1_o211440

MACRO fake_macro_adaptec1_o211441
    CLASS BLOCK ;
    SIZE 11.2 BY 299.04 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.245 0.595 294.315 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.325 0.595 290.395 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.405 0.595 286.475 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 284.165 0.595 284.235 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 280.245 0.595 280.315 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.325 0.595 276.395 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 270.725 0.595 270.795 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 266.805 0.595 266.875 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 262.885 0.595 262.955 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.645 0.595 260.715 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.725 0.595 256.795 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.805 0.595 252.875 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.205 0.595 247.275 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.285 0.595 243.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.365 0.595 239.435 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.445 0.595 235.515 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 233.205 0.595 233.275 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.285 0.595 229.355 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.685 0.595 223.755 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 219.765 0.595 219.835 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 215.845 0.595 215.915 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 211.925 0.595 211.995 ;
        END
    END p21
    PIN p22
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.685 0.595 209.755 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.765 0.595 205.835 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.845 0.595 201.915 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.245 0.595 196.315 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.325 0.595 192.395 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.405 0.595 188.475 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 186.165 0.595 186.235 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 182.245 0.595 182.315 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.325 0.595 178.395 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.405 0.595 174.475 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 168.805 0.595 168.875 ;
        END
    END p32
    PIN p33
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 164.885 0.595 164.955 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 160.965 0.595 161.035 ;
        END
    END p34
    PIN p35
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.725 0.595 158.795 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 141.085 0.595 141.155 ;
        END
    END p36
    PIN p37
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.205 0.595 135.275 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.285 0.595 131.355 ;
        END
    END p38
    PIN p39
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.365 0.595 127.435 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.405 0.595 125.475 ;
        END
    END p40
    PIN p41
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.485 0.595 121.555 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.565 0.595 117.635 ;
        END
    END p42
    PIN p43
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.645 0.595 113.715 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.765 0.595 107.835 ;
        END
    END p44
    PIN p45
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.845 0.595 103.915 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.925 0.595 99.995 ;
        END
    END p46
    PIN p47
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.965 0.595 98.035 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 94.045 0.595 94.115 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 90.125 0.595 90.195 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.245 0.595 84.315 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.325 0.595 80.395 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.405 0.595 76.475 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.485 0.595 72.555 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.525 0.595 70.595 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 60.725 0.595 60.795 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 56.805 0.595 56.875 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 52.885 0.595 52.955 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.925 0.595 50.995 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 47.005 0.595 47.075 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 43.085 0.595 43.155 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 39.165 0.595 39.235 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.285 0.595 33.355 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.365 0.595 29.435 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.445 0.595 25.515 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.485 0.595 23.555 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.565 0.595 19.635 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.645 0.595 15.715 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 9.765 0.595 9.835 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 5.845 0.595 5.915 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 1.925 0.595 1.995 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 294.525 0.595 294.595 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 153.965 9.555 154.035 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 153.685 9.555 153.755 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 152.005 9.555 152.075 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.725 0.595 151.795 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 151.165 0.595 151.235 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.645 0.595 267.715 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.565 0.595 271.635 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 275.485 0.595 275.555 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.405 0.595 279.475 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.325 0.595 283.395 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.245 0.595 287.315 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.165 0.595 291.235 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.085 0.595 295.155 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.325 0.595 143.395 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 142.205 9.555 142.275 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 169.925 9.555 169.995 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.765 0.595 2.835 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.685 0.595 6.755 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.605 0.595 10.675 ;
        END
    END p91
    PIN p92
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 14.525 0.595 14.595 ;
        END
    END p92
    PIN p93
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 18.445 0.595 18.515 ;
        END
    END p93
    PIN p94
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 22.365 0.595 22.435 ;
        END
    END p94
    PIN p95
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 26.285 0.595 26.355 ;
        END
    END p95
    PIN p96
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 30.205 0.595 30.275 ;
        END
    END p96
    PIN p97
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.125 0.595 34.195 ;
        END
    END p97
    PIN p98
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.045 0.595 38.115 ;
        END
    END p98
    PIN p99
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.965 0.595 42.035 ;
        END
    END p99
    PIN p100
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.885 0.595 45.955 ;
        END
    END p100
    PIN p101
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.805 0.595 49.875 ;
        END
    END p101
    PIN p102
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.725 0.595 53.795 ;
        END
    END p102
    PIN p103
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.645 0.595 57.715 ;
        END
    END p103
    PIN p104
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.565 0.595 61.635 ;
        END
    END p104
    PIN p105
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.485 0.595 65.555 ;
        END
    END p105
    PIN p106
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.405 0.595 69.475 ;
        END
    END p106
    PIN p107
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.325 0.595 73.395 ;
        END
    END p107
    PIN p108
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.245 0.595 77.315 ;
        END
    END p108
    PIN p109
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p109
    PIN p110
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.085 0.595 85.155 ;
        END
    END p110
    PIN p111
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p111
    PIN p112
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.925 0.595 92.995 ;
        END
    END p112
    PIN p113
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p113
    PIN p114
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.765 0.595 100.835 ;
        END
    END p114
    PIN p115
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p115
    PIN p116
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.605 0.595 108.675 ;
        END
    END p116
    PIN p117
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p117
    PIN p118
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 116.445 0.595 116.515 ;
        END
    END p118
    PIN p119
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p119
    PIN p120
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 124.285 0.595 124.355 ;
        END
    END p120
    PIN p121
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p121
    PIN p122
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.125 0.595 132.195 ;
        END
    END p122
    PIN p123
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p123
    PIN p124
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.965 0.595 140.035 ;
        END
    END p124
    PIN p125
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.885 0.595 157.955 ;
        END
    END p125
    PIN p126
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.805 0.595 161.875 ;
        END
    END p126
    PIN p127
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.725 0.595 165.795 ;
        END
    END p127
    PIN p128
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.645 0.595 169.715 ;
        END
    END p128
    PIN p129
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.565 0.595 173.635 ;
        END
    END p129
    PIN p130
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 177.485 0.595 177.555 ;
        END
    END p130
    PIN p131
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.405 0.595 181.475 ;
        END
    END p131
    PIN p132
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.325 0.595 185.395 ;
        END
    END p132
    PIN p133
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.245 0.595 189.315 ;
        END
    END p133
    PIN p134
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.165 0.595 193.235 ;
        END
    END p134
    PIN p135
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.085 0.595 197.155 ;
        END
    END p135
    PIN p136
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.005 0.595 201.075 ;
        END
    END p136
    PIN p137
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.925 0.595 204.995 ;
        END
    END p137
    PIN p138
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.845 0.595 208.915 ;
        END
    END p138
    PIN p139
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.765 0.595 212.835 ;
        END
    END p139
    PIN p140
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.685 0.595 216.755 ;
        END
    END p140
    PIN p141
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.605 0.595 220.675 ;
        END
    END p141
    PIN p142
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 224.525 0.595 224.595 ;
        END
    END p142
    PIN p143
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 228.445 0.595 228.515 ;
        END
    END p143
    PIN p144
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.365 0.595 232.435 ;
        END
    END p144
    PIN p145
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.285 0.595 236.355 ;
        END
    END p145
    PIN p146
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.205 0.595 240.275 ;
        END
    END p146
    PIN p147
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.125 0.595 244.195 ;
        END
    END p147
    PIN p148
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.045 0.595 248.115 ;
        END
    END p148
    PIN p149
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.965 0.595 252.035 ;
        END
    END p149
    PIN p150
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.885 0.595 255.955 ;
        END
    END p150
    PIN p151
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.805 0.595 259.875 ;
        END
    END p151
    PIN p152
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.725 0.595 263.795 ;
        END
    END p152
    PIN p153
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 154.245 10.115 154.315 ;
        END
    END p153
    PIN p154
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 154.805 0.595 154.875 ;
        END
    END p154
    PIN p155
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 6.125 0.595 6.195 ;
        END
    END p155
    PIN p156
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p156
    PIN p157
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p157
    PIN p158
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p158
    PIN p159
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 13.965 0.595 14.035 ;
        END
    END p159
    PIN p160
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p160
    PIN p161
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p161
    PIN p162
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p162
    PIN p163
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 21.805 0.595 21.875 ;
        END
    END p163
    PIN p164
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p164
    PIN p165
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p165
    PIN p166
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p166
    PIN p167
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 29.645 0.595 29.715 ;
        END
    END p167
    PIN p168
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p168
    PIN p169
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p169
    PIN p170
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p170
    PIN p171
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 37.485 0.595 37.555 ;
        END
    END p171
    PIN p172
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p172
    PIN p173
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p173
    PIN p174
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p174
    PIN p175
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 45.325 0.595 45.395 ;
        END
    END p175
    PIN p176
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p176
    PIN p177
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p177
    PIN p178
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p178
    PIN p179
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 53.165 0.595 53.235 ;
        END
    END p179
    PIN p180
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p180
    PIN p181
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p181
    PIN p182
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p182
    PIN p183
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 61.005 0.595 61.075 ;
        END
    END p183
    PIN p184
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p184
    PIN p185
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.925 0.595 64.995 ;
        END
    END p185
    PIN p186
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p186
    PIN p187
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.845 0.595 68.915 ;
        END
    END p187
    PIN p188
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p188
    PIN p189
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 72.765 0.595 72.835 ;
        END
    END p189
    PIN p190
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 70.245 0.595 70.315 ;
        END
    END p190
    PIN p191
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 76.685 0.595 76.755 ;
        END
    END p191
    PIN p192
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 74.165 0.595 74.235 ;
        END
    END p192
    PIN p193
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 80.605 0.595 80.675 ;
        END
    END p193
    PIN p194
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.085 0.595 78.155 ;
        END
    END p194
    PIN p195
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 84.525 0.595 84.595 ;
        END
    END p195
    PIN p196
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 82.005 0.595 82.075 ;
        END
    END p196
    PIN p197
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 88.445 0.595 88.515 ;
        END
    END p197
    PIN p198
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 85.925 0.595 85.995 ;
        END
    END p198
    PIN p199
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 92.365 0.595 92.435 ;
        END
    END p199
    PIN p200
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.845 0.595 89.915 ;
        END
    END p200
    PIN p201
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.285 0.595 96.355 ;
        END
    END p201
    PIN p202
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 93.765 0.595 93.835 ;
        END
    END p202
    PIN p203
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 100.205 0.595 100.275 ;
        END
    END p203
    PIN p204
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 97.685 0.595 97.755 ;
        END
    END p204
    PIN p205
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.125 0.595 104.195 ;
        END
    END p205
    PIN p206
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 101.605 0.595 101.675 ;
        END
    END p206
    PIN p207
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 108.045 0.595 108.115 ;
        END
    END p207
    PIN p208
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 105.525 0.595 105.595 ;
        END
    END p208
    PIN p209
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.965 0.595 112.035 ;
        END
    END p209
    PIN p210
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 109.445 0.595 109.515 ;
        END
    END p210
    PIN p211
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.885 0.595 115.955 ;
        END
    END p211
    PIN p212
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 113.365 0.595 113.435 ;
        END
    END p212
    PIN p213
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 119.805 0.595 119.875 ;
        END
    END p213
    PIN p214
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 117.285 0.595 117.355 ;
        END
    END p214
    PIN p215
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 123.725 0.595 123.795 ;
        END
    END p215
    PIN p216
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 121.205 0.595 121.275 ;
        END
    END p216
    PIN p217
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 127.645 0.595 127.715 ;
        END
    END p217
    PIN p218
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 125.125 0.595 125.195 ;
        END
    END p218
    PIN p219
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 131.565 0.595 131.635 ;
        END
    END p219
    PIN p220
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 129.045 0.595 129.115 ;
        END
    END p220
    PIN p221
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 135.485 0.595 135.555 ;
        END
    END p221
    PIN p222
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 132.965 0.595 133.035 ;
        END
    END p222
    PIN p223
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 139.405 0.595 139.475 ;
        END
    END p223
    PIN p224
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.885 0.595 136.955 ;
        END
    END p224
    PIN p225
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 158.445 0.595 158.515 ;
        END
    END p225
    PIN p226
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 140.805 0.595 140.875 ;
        END
    END p226
    PIN p227
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 162.365 0.595 162.435 ;
        END
    END p227
    PIN p228
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 157.325 0.595 157.395 ;
        END
    END p228
    PIN p229
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 166.285 0.595 166.355 ;
        END
    END p229
    PIN p230
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 161.245 0.595 161.315 ;
        END
    END p230
    PIN p231
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 170.205 0.595 170.275 ;
        END
    END p231
    PIN p232
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 165.165 0.595 165.235 ;
        END
    END p232
    PIN p233
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 174.125 0.595 174.195 ;
        END
    END p233
    PIN p234
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 169.085 0.595 169.155 ;
        END
    END p234
    PIN p235
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 178.045 0.595 178.115 ;
        END
    END p235
    PIN p236
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 173.005 0.595 173.075 ;
        END
    END p236
    PIN p237
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 181.965 0.595 182.035 ;
        END
    END p237
    PIN p238
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 176.925 0.595 176.995 ;
        END
    END p238
    PIN p239
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 185.885 0.595 185.955 ;
        END
    END p239
    PIN p240
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 180.845 0.595 180.915 ;
        END
    END p240
    PIN p241
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 189.805 0.595 189.875 ;
        END
    END p241
    PIN p242
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 184.765 0.595 184.835 ;
        END
    END p242
    PIN p243
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 193.725 0.595 193.795 ;
        END
    END p243
    PIN p244
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 188.685 0.595 188.755 ;
        END
    END p244
    PIN p245
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 197.645 0.595 197.715 ;
        END
    END p245
    PIN p246
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 192.605 0.595 192.675 ;
        END
    END p246
    PIN p247
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 201.565 0.595 201.635 ;
        END
    END p247
    PIN p248
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 196.525 0.595 196.595 ;
        END
    END p248
    PIN p249
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 205.485 0.595 205.555 ;
        END
    END p249
    PIN p250
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 200.445 0.595 200.515 ;
        END
    END p250
    PIN p251
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 209.405 0.595 209.475 ;
        END
    END p251
    PIN p252
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 204.365 0.595 204.435 ;
        END
    END p252
    PIN p253
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 213.325 0.595 213.395 ;
        END
    END p253
    PIN p254
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 208.285 0.595 208.355 ;
        END
    END p254
    PIN p255
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 217.245 0.595 217.315 ;
        END
    END p255
    PIN p256
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 212.205 0.595 212.275 ;
        END
    END p256
    PIN p257
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 221.165 0.595 221.235 ;
        END
    END p257
    PIN p258
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 216.125 0.595 216.195 ;
        END
    END p258
    PIN p259
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 225.085 0.595 225.155 ;
        END
    END p259
    PIN p260
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 220.045 0.595 220.115 ;
        END
    END p260
    PIN p261
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 229.005 0.595 229.075 ;
        END
    END p261
    PIN p262
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 223.965 0.595 224.035 ;
        END
    END p262
    PIN p263
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 232.925 0.595 232.995 ;
        END
    END p263
    PIN p264
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 227.885 0.595 227.955 ;
        END
    END p264
    PIN p265
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 236.845 0.595 236.915 ;
        END
    END p265
    PIN p266
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 231.805 0.595 231.875 ;
        END
    END p266
    PIN p267
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 240.765 0.595 240.835 ;
        END
    END p267
    PIN p268
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 235.725 0.595 235.795 ;
        END
    END p268
    PIN p269
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 244.685 0.595 244.755 ;
        END
    END p269
    PIN p270
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 239.645 0.595 239.715 ;
        END
    END p270
    PIN p271
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 248.605 0.595 248.675 ;
        END
    END p271
    PIN p272
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 243.565 0.595 243.635 ;
        END
    END p272
    PIN p273
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 252.525 0.595 252.595 ;
        END
    END p273
    PIN p274
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 247.485 0.595 247.555 ;
        END
    END p274
    PIN p275
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 256.445 0.595 256.515 ;
        END
    END p275
    PIN p276
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 251.405 0.595 251.475 ;
        END
    END p276
    PIN p277
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 260.365 0.595 260.435 ;
        END
    END p277
    PIN p278
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 255.325 0.595 255.395 ;
        END
    END p278
    PIN p279
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 264.285 0.595 264.355 ;
        END
    END p279
    PIN p280
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 259.245 0.595 259.315 ;
        END
    END p280
    PIN p281
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 268.205 0.595 268.275 ;
        END
    END p281
    PIN p282
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 263.165 0.595 263.235 ;
        END
    END p282
    PIN p283
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 272.125 0.595 272.195 ;
        END
    END p283
    PIN p284
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 267.085 0.595 267.155 ;
        END
    END p284
    PIN p285
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 276.045 0.595 276.115 ;
        END
    END p285
    PIN p286
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 271.005 0.595 271.075 ;
        END
    END p286
    PIN p287
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 279.965 0.595 280.035 ;
        END
    END p287
    PIN p288
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 274.925 0.595 274.995 ;
        END
    END p288
    PIN p289
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 283.885 0.595 283.955 ;
        END
    END p289
    PIN p290
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 278.845 0.595 278.915 ;
        END
    END p290
    PIN p291
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 287.805 0.595 287.875 ;
        END
    END p291
    PIN p292
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 282.765 0.595 282.835 ;
        END
    END p292
    PIN p293
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 291.725 0.595 291.795 ;
        END
    END p293
    PIN p294
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 286.685 0.595 286.755 ;
        END
    END p294
    PIN p295
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 295.645 0.595 295.715 ;
        END
    END p295
    PIN p296
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 290.605 0.595 290.675 ;
        END
    END p296
    PIN p297
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 85.085 9.555 85.155 ;
        END
    END p297
    PIN p298
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 81.165 9.555 81.235 ;
        END
    END p298
    PIN p299
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 77.245 9.555 77.315 ;
        END
    END p299
    PIN p300
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 73.325 9.555 73.395 ;
        END
    END p300
    PIN p301
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 69.405 9.555 69.475 ;
        END
    END p301
    PIN p302
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 65.485 9.555 65.555 ;
        END
    END p302
    PIN p303
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 61.565 9.555 61.635 ;
        END
    END p303
    PIN p304
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 57.645 9.555 57.715 ;
        END
    END p304
    PIN p305
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 53.725 9.555 53.795 ;
        END
    END p305
    PIN p306
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 49.805 9.555 49.875 ;
        END
    END p306
    PIN p307
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 45.885 9.555 45.955 ;
        END
    END p307
    PIN p308
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 41.965 9.555 42.035 ;
        END
    END p308
    PIN p309
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 38.045 9.555 38.115 ;
        END
    END p309
    PIN p310
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 34.125 9.555 34.195 ;
        END
    END p310
    PIN p311
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 30.205 9.555 30.275 ;
        END
    END p311
    PIN p312
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 26.285 9.555 26.355 ;
        END
    END p312
    PIN p313
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 22.365 9.555 22.435 ;
        END
    END p313
    PIN p314
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 18.445 9.555 18.515 ;
        END
    END p314
    PIN p315
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 14.525 9.555 14.595 ;
        END
    END p315
    PIN p316
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 10.605 9.555 10.675 ;
        END
    END p316
    PIN p317
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 6.685 9.555 6.755 ;
        END
    END p317
    PIN p318
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 2.765 9.555 2.835 ;
        END
    END p318
    PIN p319
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 255.885 9.555 255.955 ;
        END
    END p319
    PIN p320
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 251.965 9.555 252.035 ;
        END
    END p320
    PIN p321
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 248.045 9.555 248.115 ;
        END
    END p321
    PIN p322
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 244.125 9.555 244.195 ;
        END
    END p322
    PIN p323
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 240.205 9.555 240.275 ;
        END
    END p323
    PIN p324
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 236.285 9.555 236.355 ;
        END
    END p324
    PIN p325
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 232.365 9.555 232.435 ;
        END
    END p325
    PIN p326
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 228.445 9.555 228.515 ;
        END
    END p326
    PIN p327
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 224.525 9.555 224.595 ;
        END
    END p327
    PIN p328
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 220.605 9.555 220.675 ;
        END
    END p328
    PIN p329
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 216.685 9.555 216.755 ;
        END
    END p329
    PIN p330
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 212.765 9.555 212.835 ;
        END
    END p330
    PIN p331
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 208.845 9.555 208.915 ;
        END
    END p331
    PIN p332
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 204.925 9.555 204.995 ;
        END
    END p332
    PIN p333
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 201.005 9.555 201.075 ;
        END
    END p333
    PIN p334
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 197.085 9.555 197.155 ;
        END
    END p334
    PIN p335
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 193.165 9.555 193.235 ;
        END
    END p335
    PIN p336
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 189.245 9.555 189.315 ;
        END
    END p336
    PIN p337
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 185.325 9.555 185.395 ;
        END
    END p337
    PIN p338
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 181.405 9.555 181.475 ;
        END
    END p338
    PIN p339
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 295.085 9.555 295.155 ;
        END
    END p339
    PIN p340
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 291.165 9.555 291.235 ;
        END
    END p340
    PIN p341
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 287.245 9.555 287.315 ;
        END
    END p341
    PIN p342
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 283.325 9.555 283.395 ;
        END
    END p342
    PIN p343
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 279.405 9.555 279.475 ;
        END
    END p343
    PIN p344
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 275.485 9.555 275.555 ;
        END
    END p344
    PIN p345
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 271.565 9.555 271.635 ;
        END
    END p345
    PIN p346
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 177.485 9.555 177.555 ;
        END
    END p346
    PIN p347
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 267.645 9.555 267.715 ;
        END
    END p347
    PIN p348
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 173.565 9.555 173.635 ;
        END
    END p348
    PIN p349
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 263.725 9.555 263.795 ;
        END
    END p349
    PIN p350
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 169.645 9.555 169.715 ;
        END
    END p350
    PIN p351
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 259.805 9.555 259.875 ;
        END
    END p351
    PIN p352
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 165.725 9.555 165.795 ;
        END
    END p352
    PIN p353
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 161.805 9.555 161.875 ;
        END
    END p353
    PIN p354
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 157.885 9.555 157.955 ;
        END
    END p354
    PIN p355
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 139.965 9.555 140.035 ;
        END
    END p355
    PIN p356
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 136.045 9.555 136.115 ;
        END
    END p356
    PIN p357
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 132.125 9.555 132.195 ;
        END
    END p357
    PIN p358
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 128.205 9.555 128.275 ;
        END
    END p358
    PIN p359
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 124.285 9.555 124.355 ;
        END
    END p359
    PIN p360
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 120.365 9.555 120.435 ;
        END
    END p360
    PIN p361
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 116.445 9.555 116.515 ;
        END
    END p361
    PIN p362
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 112.525 9.555 112.595 ;
        END
    END p362
    PIN p363
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 108.605 9.555 108.675 ;
        END
    END p363
    PIN p364
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 104.685 9.555 104.755 ;
        END
    END p364
    PIN p365
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 100.765 9.555 100.835 ;
        END
    END p365
    PIN p366
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 96.845 9.555 96.915 ;
        END
    END p366
    PIN p367
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 92.925 9.555 92.995 ;
        END
    END p367
    PIN p368
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  9.485 89.005 9.555 89.075 ;
        END
    END p368
    PIN p369
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p369
    OBS
      LAYER via2 ;
        RECT  0 0 11.2 299.04 ;
      LAYER metal2 ;
        RECT  0 0 11.2 299.04 ;
      LAYER via1 ;
        RECT  0 0 11.2 299.04 ;
      LAYER metal1 ;
        RECT  0 0 11.2 299.04 ;
    END
END fake_macro_adaptec1_o211441

MACRO fake_macro_adaptec1_o211442
    CLASS BLOCK ;
    SIZE 100.8 BY 147.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 138.005 2.275 138.075 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 130.165 2.275 130.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 122.325 2.275 122.395 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 114.485 2.275 114.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 106.645 2.275 106.715 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 98.805 2.275 98.875 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 90.965 2.275 91.035 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 83.125 2.275 83.195 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 79.765 96.355 79.835 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.885 0.595 143.955 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.045 0.595 115.115 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.525 0.595 91.595 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p27
    PIN p28
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p29
    PIN p30
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.685 0.595 83.755 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.365 0.595 99.435 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.205 0.595 107.275 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.885 0.595 122.955 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.725 0.595 130.795 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.565 0.595 138.635 ;
        END
    END p48
    PIN p49
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 76.405 96.915 76.475 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 69.965 96.915 70.035 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.885 0.595 66.955 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 67.725 0.595 67.795 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.965 0.595 70.035 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.005 0.595 68.075 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.725 0.595 95.795 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 67.445 0.595 67.515 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 78.645 97.475 78.715 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 73.885 97.475 73.955 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.805 0.595 77.875 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.605 0.595 73.675 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.445 0.595 81.515 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.885 0.595 73.955 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.885 1.155 73.955 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 80.605 96.355 80.675 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.365 0.595 64.435 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.765 0.595 65.835 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 64.085 96.355 64.155 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 63.805 96.355 63.875 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 67.165 1.155 67.235 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.605 0.595 87.675 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.445 0.595 95.515 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.285 0.595 103.355 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.125 0.595 111.195 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.965 0.595 119.035 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.805 0.595 126.875 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.645 0.595 134.715 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.485 0.595 142.555 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 108.325 96.355 108.395 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 6.685 98.595 6.755 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 14.525 98.595 14.595 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 22.365 98.595 22.435 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 30.205 98.595 30.275 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 38.045 98.595 38.115 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 6.125 99.155 6.195 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 45.885 98.595 45.955 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 13.965 99.155 14.035 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 53.725 98.595 53.795 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 21.805 99.155 21.875 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 61.565 98.595 61.635 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 29.645 99.155 29.715 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 84.525 98.595 84.595 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 37.485 99.155 37.555 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 92.365 98.595 92.435 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 45.325 99.155 45.395 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 53.165 99.155 53.235 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 61.005 99.155 61.075 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 85.085 99.155 85.155 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 92.925 99.155 92.995 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 100.765 99.155 100.835 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 108.605 99.155 108.675 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 116.445 99.155 116.515 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 124.285 99.155 124.355 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 132.125 99.155 132.195 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 139.965 99.155 140.035 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 100.205 98.595 100.275 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 108.045 98.595 108.115 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 115.885 98.595 115.955 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 123.725 98.595 123.795 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 131.565 98.595 131.635 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 139.405 98.595 139.475 ;
        END
    END p123
    OBS
      LAYER via2 ;
        RECT  0 0 100.8 147.84 ;
      LAYER metal2 ;
        RECT  0 0 100.8 147.84 ;
      LAYER via1 ;
        RECT  0 0 100.8 147.84 ;
      LAYER metal1 ;
        RECT  0 0 100.8 147.84 ;
    END
END fake_macro_adaptec1_o211442

MACRO fake_macro_adaptec1_o211443
    CLASS BLOCK ;
    SIZE 100.8 BY 147.84 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 138.005 2.275 138.075 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 130.165 2.275 130.235 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 122.325 2.275 122.395 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 114.485 2.275 114.555 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 106.645 2.275 106.715 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 98.805 2.275 98.875 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 90.965 2.275 91.035 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 83.125 2.275 83.195 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 56.525 2.275 56.595 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 48.685 2.275 48.755 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 40.845 2.275 40.915 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 33.005 2.275 33.075 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 25.165 2.275 25.235 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 17.325 2.275 17.395 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 9.485 2.275 9.555 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  2.205 1.645 2.275 1.715 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 79.765 96.355 79.835 ;
        END
    END p16
    PIN p17
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 41.405 0.595 41.475 ;
        END
    END p17
    PIN p18
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 17.885 0.595 17.955 ;
        END
    END p18
    PIN p19
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 143.885 0.595 143.955 ;
        END
    END p19
    PIN p20
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 89.005 0.595 89.075 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 7.525 0.595 7.595 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 112.525 0.595 112.595 ;
        END
    END p22
    PIN p23
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 115.045 0.595 115.115 ;
        END
    END p23
    PIN p24
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 91.525 0.595 91.595 ;
        END
    END p24
    PIN p25
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 54.565 0.595 54.635 ;
        END
    END p25
    PIN p26
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 80.605 96.355 80.675 ;
        END
    END p26
    PIN p27
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 108.325 96.355 108.395 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 2.205 0.595 2.275 ;
        END
    END p28
    PIN p29
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 15.365 0.595 15.435 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 10.045 0.595 10.115 ;
        END
    END p30
    PIN p31
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 23.205 0.595 23.275 ;
        END
    END p31
    PIN p32
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 31.045 0.595 31.115 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 25.725 0.595 25.795 ;
        END
    END p33
    PIN p34
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 38.885 0.595 38.955 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 33.565 0.595 33.635 ;
        END
    END p35
    PIN p36
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 46.725 0.595 46.795 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 49.245 0.595 49.315 ;
        END
    END p37
    PIN p38
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 62.405 0.595 62.475 ;
        END
    END p38
    PIN p39
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 57.085 0.595 57.155 ;
        END
    END p39
    PIN p40
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 83.685 0.595 83.755 ;
        END
    END p40
    PIN p41
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 96.845 0.595 96.915 ;
        END
    END p41
    PIN p42
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 99.365 0.595 99.435 ;
        END
    END p42
    PIN p43
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 104.685 0.595 104.755 ;
        END
    END p43
    PIN p44
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 107.205 0.595 107.275 ;
        END
    END p44
    PIN p45
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 120.365 0.595 120.435 ;
        END
    END p45
    PIN p46
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 122.885 0.595 122.955 ;
        END
    END p46
    PIN p47
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 128.205 0.595 128.275 ;
        END
    END p47
    PIN p48
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 130.725 0.595 130.795 ;
        END
    END p48
    PIN p49
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 136.045 0.595 136.115 ;
        END
    END p49
    PIN p50
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 138.565 0.595 138.635 ;
        END
    END p50
    PIN p51
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 76.405 96.915 76.475 ;
        END
    END p51
    PIN p52
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.845 69.965 96.915 70.035 ;
        END
    END p52
    PIN p53
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.885 0.595 66.955 ;
        END
    END p53
    PIN p54
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 67.725 0.595 67.795 ;
        END
    END p54
    PIN p55
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 69.965 0.595 70.035 ;
        END
    END p55
    PIN p56
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 68.005 0.595 68.075 ;
        END
    END p56
    PIN p57
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.725 0.595 95.795 ;
        END
    END p57
    PIN p58
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 67.445 0.595 67.515 ;
        END
    END p58
    PIN p59
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 78.645 97.475 78.715 ;
        END
    END p59
    PIN p60
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  97.405 73.885 97.475 73.955 ;
        END
    END p60
    PIN p61
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 78.365 0.595 78.435 ;
        END
    END p61
    PIN p62
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 77.805 0.595 77.875 ;
        END
    END p62
    PIN p63
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.605 0.595 73.675 ;
        END
    END p63
    PIN p64
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.445 0.595 81.515 ;
        END
    END p64
    PIN p65
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 73.885 0.595 73.955 ;
        END
    END p65
    PIN p66
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 73.885 1.155 73.955 ;
        END
    END p66
    PIN p67
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 64.365 0.595 64.435 ;
        END
    END p67
    PIN p68
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 65.765 0.595 65.835 ;
        END
    END p68
    PIN p69
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 64.085 96.355 64.155 ;
        END
    END p69
    PIN p70
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  96.285 63.805 96.355 63.875 ;
        END
    END p70
    PIN p71
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.325 0.595 66.395 ;
        END
    END p71
    PIN p72
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 67.165 1.155 67.235 ;
        END
    END p72
    PIN p73
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 66.605 0.595 66.675 ;
        END
    END p73
    PIN p74
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  1.085 66.885 1.155 66.955 ;
        END
    END p74
    PIN p75
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 3.605 0.595 3.675 ;
        END
    END p75
    PIN p76
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 11.445 0.595 11.515 ;
        END
    END p76
    PIN p77
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 19.285 0.595 19.355 ;
        END
    END p77
    PIN p78
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 27.125 0.595 27.195 ;
        END
    END p78
    PIN p79
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 34.965 0.595 35.035 ;
        END
    END p79
    PIN p80
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 42.805 0.595 42.875 ;
        END
    END p80
    PIN p81
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 50.645 0.595 50.715 ;
        END
    END p81
    PIN p82
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 58.485 0.595 58.555 ;
        END
    END p82
    PIN p83
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 87.605 0.595 87.675 ;
        END
    END p83
    PIN p84
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 95.445 0.595 95.515 ;
        END
    END p84
    PIN p85
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 103.285 0.595 103.355 ;
        END
    END p85
    PIN p86
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 111.125 0.595 111.195 ;
        END
    END p86
    PIN p87
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 118.965 0.595 119.035 ;
        END
    END p87
    PIN p88
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 126.805 0.595 126.875 ;
        END
    END p88
    PIN p89
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 134.645 0.595 134.715 ;
        END
    END p89
    PIN p90
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 142.485 0.595 142.555 ;
        END
    END p90
    PIN p91
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  0.525 81.165 0.595 81.235 ;
        END
    END p91
    PIN p92
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 6.685 98.595 6.755 ;
        END
    END p92
    PIN p93
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 14.525 98.595 14.595 ;
        END
    END p93
    PIN p94
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 22.365 98.595 22.435 ;
        END
    END p94
    PIN p95
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 30.205 98.595 30.275 ;
        END
    END p95
    PIN p96
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 38.045 98.595 38.115 ;
        END
    END p96
    PIN p97
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 6.125 99.155 6.195 ;
        END
    END p97
    PIN p98
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 45.885 98.595 45.955 ;
        END
    END p98
    PIN p99
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 13.965 99.155 14.035 ;
        END
    END p99
    PIN p100
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 53.725 98.595 53.795 ;
        END
    END p100
    PIN p101
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 21.805 99.155 21.875 ;
        END
    END p101
    PIN p102
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 61.565 98.595 61.635 ;
        END
    END p102
    PIN p103
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 29.645 99.155 29.715 ;
        END
    END p103
    PIN p104
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 84.525 98.595 84.595 ;
        END
    END p104
    PIN p105
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 37.485 99.155 37.555 ;
        END
    END p105
    PIN p106
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 92.365 98.595 92.435 ;
        END
    END p106
    PIN p107
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 45.325 99.155 45.395 ;
        END
    END p107
    PIN p108
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 53.165 99.155 53.235 ;
        END
    END p108
    PIN p109
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 61.005 99.155 61.075 ;
        END
    END p109
    PIN p110
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 85.085 99.155 85.155 ;
        END
    END p110
    PIN p111
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 92.925 99.155 92.995 ;
        END
    END p111
    PIN p112
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 100.765 99.155 100.835 ;
        END
    END p112
    PIN p113
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 108.605 99.155 108.675 ;
        END
    END p113
    PIN p114
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 116.445 99.155 116.515 ;
        END
    END p114
    PIN p115
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 124.285 99.155 124.355 ;
        END
    END p115
    PIN p116
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 132.125 99.155 132.195 ;
        END
    END p116
    PIN p117
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  99.085 139.965 99.155 140.035 ;
        END
    END p117
    PIN p118
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 100.205 98.595 100.275 ;
        END
    END p118
    PIN p119
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 108.045 98.595 108.115 ;
        END
    END p119
    PIN p120
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 115.885 98.595 115.955 ;
        END
    END p120
    PIN p121
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 123.725 98.595 123.795 ;
        END
    END p121
    PIN p122
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 131.565 98.595 131.635 ;
        END
    END p122
    PIN p123
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  98.525 139.405 98.595 139.475 ;
        END
    END p123
    OBS
      LAYER via2 ;
        RECT  0 0 100.8 147.84 ;
      LAYER metal2 ;
        RECT  0 0 100.8 147.84 ;
      LAYER via1 ;
        RECT  0 0 100.8 147.84 ;
      LAYER metal1 ;
        RECT  0 0 100.8 147.84 ;
    END
END fake_macro_adaptec1_o211443

MACRO fake_macro_adaptec1_o211444
    CLASS BLOCK ;
    SIZE 146.72 BY 114.24 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 107.765 81.795 107.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 107.765 75.635 107.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.805 107.765 77.875 107.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.885 107.765 73.955 107.835 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 107.765 82.355 107.835 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.165 107.765 81.235 107.835 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 107.765 71.715 107.835 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.205 107.765 72.275 107.835 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 107.765 73.395 107.835 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 12.285 10.115 12.355 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  74.445 6.125 74.515 6.195 ;
        END
    END p10
    PIN p11
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 107.765 66.675 107.835 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 107.765 64.995 107.835 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.245 107.765 77.315 107.835 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 107.765 79.555 107.835 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.125 107.765 76.195 107.835 ;
        END
    END p15
    PIN p16
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 107.765 78.995 107.835 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 107.765 67.235 107.835 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.045 107.765 80.115 107.835 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 107.765 80.675 107.835 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 113.925 80.675 113.995 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 107.765 63.875 107.835 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.365 107.765 78.435 107.835 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 113.925 78.995 113.995 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 113.925 64.995 113.995 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 107.485 67.795 107.555 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  134.365 107.485 134.435 107.555 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 107.765 64.435 107.835 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.085 107.765 71.155 107.835 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.205 113.925 72.275 113.995 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.765 107.765 72.835 107.835 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.885 113.925 73.955 113.995 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 107.765 75.075 107.835 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.565 113.925 75.635 113.995 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  76.685 107.765 76.755 107.835 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  77.245 113.925 77.315 113.995 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 107.765 65.555 107.835 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  125.965 107.765 126.035 107.835 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  10.045 107.485 10.115 107.555 ;
        END
    END p38
    OBS
      LAYER via2 ;
        RECT  0 0 146.72 114.24 ;
      LAYER metal2 ;
        RECT  0 0 146.72 114.24 ;
      LAYER via1 ;
        RECT  0 0 146.72 114.24 ;
      LAYER metal1 ;
        RECT  0 0 146.72 114.24 ;
    END
END fake_macro_adaptec1_o211444

MACRO fake_macro_adaptec1_o211445
    CLASS BLOCK ;
    SIZE 146.72 BY 114.24 ;
    SYMMETRY X Y ;
    PIN p0
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.365 107.765 64.435 107.835 ;
        END
    END p0
    PIN p1
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 107.765 70.595 107.835 ;
        END
    END p1
    PIN p2
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.965 107.765 70.035 107.835 ;
        END
    END p2
    PIN p3
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.285 107.765 68.355 107.835 ;
        END
    END p3
    PIN p4
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 107.765 67.235 107.835 ;
        END
    END p4
    PIN p5
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.205 107.765 72.275 107.835 ;
        END
    END p5
    PIN p6
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  63.805 107.765 63.875 107.835 ;
        END
    END p6
    PIN p7
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  64.925 107.765 64.995 107.835 ;
        END
    END p7
    PIN p8
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 107.765 68.915 107.835 ;
        END
    END p8
    PIN p9
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.605 107.765 66.675 107.835 ;
        END
    END p9
    PIN p10
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  74.445 107.765 74.515 107.835 ;
        END
    END p10
    PIN p11
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.885 107.765 73.955 107.835 ;
        END
    END p11
    PIN p12
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.765 107.765 72.835 107.835 ;
        END
    END p12
    PIN p13
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 12.285 136.115 12.355 ;
        END
    END p13
    PIN p14
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.645 6.125 71.715 6.195 ;
        END
    END p14
    PIN p15
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  82.285 107.765 82.355 107.835 ;
        END
    END p15
    PIN p16
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  79.485 107.765 79.555 107.835 ;
        END
    END p16
    PIN p17
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  66.045 107.765 66.115 107.835 ;
        END
    END p17
    PIN p18
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 107.765 65.555 107.835 ;
        END
    END p18
    PIN p19
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  65.485 113.925 65.555 113.995 ;
        END
    END p19
    PIN p20
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.165 107.765 81.235 107.835 ;
        END
    END p20
    PIN p21
        DIRECTION INPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.925 107.765 78.995 107.835 ;
        END
    END p21
    PIN p22
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  78.365 107.485 78.435 107.555 ;
        END
    END p22
    PIN p23
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.725 107.765 81.795 107.835 ;
        END
    END p23
    PIN p24
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  75.005 107.765 75.075 107.835 ;
        END
    END p24
    PIN p25
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.885 113.925 73.955 113.995 ;
        END
    END p25
    PIN p26
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  73.325 107.765 73.395 107.835 ;
        END
    END p26
    PIN p27
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  72.205 113.925 72.275 113.995 ;
        END
    END p27
    PIN p28
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  71.085 107.765 71.155 107.835 ;
        END
    END p28
    PIN p29
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  70.525 113.925 70.595 113.995 ;
        END
    END p29
    PIN p30
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  69.405 107.765 69.475 107.835 ;
        END
    END p30
    PIN p31
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  68.845 113.925 68.915 113.995 ;
        END
    END p31
    PIN p32
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.725 107.765 67.795 107.835 ;
        END
    END p32
    PIN p33
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  11.725 107.485 11.795 107.555 ;
        END
    END p33
    PIN p34
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  67.165 113.925 67.235 113.995 ;
        END
    END p34
    PIN p35
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  81.165 113.925 81.235 113.995 ;
        END
    END p35
    PIN p36
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  80.605 107.765 80.675 107.835 ;
        END
    END p36
    PIN p37
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  20.125 107.765 20.195 107.835 ;
        END
    END p37
    PIN p38
        DIRECTION OUTPUT ; 
        USE SIGNAL ; 
        PORT
            LAYER metal3 ;
              RECT  136.045 107.485 136.115 107.555 ;
        END
    END p38
    OBS
      LAYER via2 ;
        RECT  0 0 146.72 114.24 ;
      LAYER metal2 ;
        RECT  0 0 146.72 114.24 ;
      LAYER via1 ;
        RECT  0 0 146.72 114.24 ;
      LAYER metal1 ;
        RECT  0 0 146.72 114.24 ;
    END
END fake_macro_adaptec1_o211445
END LIBRARY
